**** Created by MC2: Version 2012.02.00.d on 2024/01/10, 17:25:26 

************************************************************************
* AUCDL NETLIST:
* 
* LIBRARY NAME:  N28HPM_DP_LEAFCELLS
* TOP CELL NAME: LEAFCELL_DP
* VIEW NAME:     SCHEMATIC
* NETLISTED ON:  DEC 24 13:14:24 2013
************************************************************************

*.EQUATION
*.SCALE METER
.PARAM


*.PIN VSS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    INV_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_INV_BULK A G GB P PB Y
*.PININFO A:I G:I GB:I P:I PB:I Y:O
M1 Y A P PB pch_mac L=LP W=WP M=MULTI*FP
M3 Y A G GB nch_mac L=LN W=WN M=MULTI*FN
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DIN_WOBIST_DP_V2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DIN_WOBIST_DP_V2 BWEB CKD D DCLKA GW GWB VDDI VSSI
*.PININFO BWEB:I CKD:I D:I DCLKA:I GW:O GWB:O VDDI:B VSSI:B
MM29 DX4L DCLKA1B Z6 VDDI pch_mac L=30N W=320N M=1
MM5 NET0129 BWEB Z13 VDDI pch_mac L=30N W=320N M=1
MM6 VDDI BX4L1B Z16 VDDI pch_mac L=30N W=320N M=1
MM27 DX4L D Z9 VDDI pch_mac L=30N W=320N M=1
MP1 DX4L3B_AND CKD2 VDDI VDDI pch_mac L=30N W=350N M=1
MM54 DX4L3B_AND BX4L1B VDDI VDDI pch_mac L=30N W=350N M=1
MM53 DX4L2_AND BX4L1B VDDI VDDI pch_mac L=30N W=350N M=1
MM52 DX4L2_AND NET108 VDDI VDDI pch_mac L=30N W=350N M=1
MM51 DX4L3B_AND DX4L2 VDDI VDDI pch_mac L=30N W=350N M=1
MM28 VDDI NET108 Z6 VDDI pch_mac L=30N W=320N M=1
MP10 DX4L2_AND CKD2 VDDI VDDI pch_mac L=30N W=350N M=1
MM7 VDDI DCLKA2 Z13 VDDI pch_mac L=30N W=320N M=1
MM4 NET0129 DCLKA1B Z16 VDDI pch_mac L=30N W=320N M=1
MM26 VDDI DCLKA2 Z9 VDDI pch_mac L=30N W=320N M=1
MM3 NET0129 BWEB Z15 VSSI nch_mac L=30N W=210N M=1
MM34 DX4L D Z11 VSSI nch_mac L=30N W=210N M=1
MM35 DX4L DCLKA2 Z7 VSSI nch_mac L=30N W=210N M=1
MM2 NET0129 DCLKA2 Z14 VSSI nch_mac L=30N W=210N M=1
MN2 Z2 CKD2 Z1 VSSI nch_mac L=30N W=760N M=2
MN33 DX4L3B_AND DX4L2 Z2 VSSI nch_mac L=30N W=760N M=1
MM1 VSSI DCLKA1B Z15 VSSI nch_mac L=30N W=210N M=1
MM37 VSSI NET108 Z7 VSSI nch_mac L=30N W=210N M=1
MM36 VSSI DCLKA1B Z11 VSSI nch_mac L=30N W=210N M=1
MM0 VSSI BX4L1B Z14 VSSI nch_mac L=30N W=210N M=1
MN1 DX4L2_AND NET108 Z2 VSSI nch_mac L=30N W=760N M=1
MN7 Z1 BX4L1B VSSI VSSI nch_mac L=30N W=1.01U M=3
XI331 NET108 VSSI VSSI VDDI VDDI DX4L2 SDBM200W80_INV_BULK FN=1 WN=0.64U LN=0.03U 
+ MULTI=1 FP=1 WP=0.98U LP=0.03U
XI314 CKD VSSI VSSI VDDI VDDI CKD1B SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI317 CKD1B VSSI VSSI VDDI VDDI CKD2 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U MULTI=1 
+ FP=1 WP=0.64U LP=0.03U
XI339 DCLKA1B VSSI VSSI VDDI VDDI DCLKA2 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U 
+ MULTI=1 FP=1 WP=0.64U LP=0.03U
XI333 DX4L3B_AND VSSI VSSI VDDI VDDI GW SDBM200W80_INV_BULK FN=10 WN=0.225U LN=0.03U 
+ MULTI=1 FP=10 WP=0.45U LP=0.03U
XI337 DCLKA VSSI VSSI VDDI VDDI DCLKA1B SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.32U LP=0.03U
XI332 DX4L2_AND VSSI VSSI VDDI VDDI GWB SDBM200W80_INV_BULK FN=10 WN=0.225U LN=0.03U 
+ MULTI=1 FP=10 WP=0.45U LP=0.03U
XI329 DX4L VSSI VSSI VDDI VDDI NET108 SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U 
+ MULTI=1 FP=1 WP=0.54U LP=0.03U
XI336 NET0129 VSSI VSSI VDDI VDDI BX4L1B SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U 
+ MULTI=1 FP=1 WP=0.54U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    NOR_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_NOR_BULK A B G GB P PB Y
*.PININFO A:I B:I G:I GB:I P:I PB:I Y:O
M1 NET021 A P PB pch_mac L=LP1 W=WP1 M=MULTI*FP1
M3 Y B NET021 PB pch_mac L=LP2 W=WP2 M=MULTI*FP2
M5 Y B G GB nch_mac L=LN2 W=WN2 M=MULTI*FN2
M7 Y A G GB nch_mac L=LN1 W=WN1 M=MULTI*FN1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DOUT_DP_V1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DOUT_DP_V1 AWT AWTDA AWTDB GBL GBLB QA QB QLATCH_AB QLATCH_BB VDDI 
+ VSSI WLP_SAEB
*.PININFO AWT:I AWTDA:I AWTDB:I QLATCH_AB:I QLATCH_BB:I WLP_SAEB:I QA:O QB:O 
*.PININFO GBL:B GBLB:B VDDI:B VSSI:B
XI216 SEL_B VSSI VSSI VDDI VDDI SEL_BB SDBM200W80_INV_BULK FN=1 WN=0.24U LN=0.03U 
+ MULTI=1 FP=2 WP=0.25U LP=0.03U
XI215 SEL_A VSSI VSSI VDDI VDDI SEL_AB SDBM200W80_INV_BULK FN=1 WN=0.24U LN=0.03U 
+ MULTI=1 FP=2 WP=0.25U LP=0.03U
XI208 QBB VSSI VSSI VDDI VDDI QBBB SDBM200W80_INV_BULK FN=1 WN=0.3U LN=0.03U MULTI=1 
+ FP=1 WP=0.4U LP=0.03U
XI205 AWTDB1B VSSI VSSI VDDI VDDI NET0173 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI200 QAB VSSI VSSI VDDI VDDI QABB SDBM200W80_INV_BULK FN=1 WN=0.3U LN=0.03U MULTI=1 
+ FP=1 WP=0.4U LP=0.03U
XI204 AWTDB VSSI VSSI VDDI VDDI AWTDB1B SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.22U LP=0.03U
XI176 SEL_A VSSI VSSI VDDI VDDI SEL_AB SDBM200W80_INV_BULK FN=1 WN=0.24U LN=0.03U 
+ MULTI=1 FP=1 WP=0.48U LP=0.03U
XI212 AWT VSSI VSSI VDDI VDDI AWT1B SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 
+ FP=1 WP=0.22U LP=0.03U
XI217 WLP_SAEB VSSI VSSI VDDI VDDI NET0229 SDBM200W80_INV_BULK FN=1 WN=0.25U LN=0.03U 
+ MULTI=1 FP=1 WP=0.25U LP=0.03U
XINV3 NET0229 VSSI VSSI VDDI VDDI DLRSB SDBM200W80_INV_BULK FN=1 WN=0.87U LN=0.03U 
+ MULTI=1 FP=1 WP=0.93U LP=0.03U
XI118 AWTDA1B VSSI VSSI VDDI VDDI NET085 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI213 AWT1B VSSI VSSI VDDI VDDI AWT2 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 
+ FP=1 WP=0.22U LP=0.03U
XI209 SEL_B VSSI VSSI VDDI VDDI SEL_BB SDBM200W80_INV_BULK FN=1 WN=0.24U LN=0.03U 
+ MULTI=1 FP=1 WP=0.48U LP=0.03U
XI207 QBB VSSI VSSI VDDI VDDI QB SDBM200W80_INV_BULK FN=4 WN=0.22U LN=0.03U MULTI=1 
+ FP=2 WP=0.8U LP=0.03U
XI198 QAB VSSI VSSI VDDI VDDI QA SDBM200W80_INV_BULK FN=4 WN=0.22U LN=0.03U MULTI=1 
+ FP=2 WP=0.8U LP=0.03U
XINV0 AWTDA VSSI VSSI VDDI VDDI AWTDA1B SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.22U LP=0.03U
MM51 NET0219 AWT1B VSSI VSSI nch_mac L=30N W=220N M=1
MM49 NET0205 AWT1B VSSI VSSI nch_mac L=30N W=220N M=1
MM40 NET0197 SEL_B VSSI VSSI nch_mac L=30N W=0.3U M=6
MM42 QBB QB_T NET0197 VSSI nch_mac L=30N W=300N M=3
MM37 QBB AWT2 NET067 VSSI nch_mac L=30N W=300N M=1
MM43 QBB QBBB NET0196 VSSI nch_mac L=30N W=220N M=1
MM31 QAB QB_T NET0145 VSSI nch_mac L=30N W=300N M=3
MM26 NET0145 SEL_A VSSI VSSI nch_mac L=30N W=0.3U M=6
MM41 NET0196 SEL_BB NET0219 VSSI nch_mac L=30N W=220N M=1
MM24 Z3 GBLB VSSI VSSI nch_mac L=30N W=0.33U M=4
MM36 NET067 NET0173 VSSI VSSI nch_mac L=30N W=300N M=1
MM32 QAB QABB NET0144 VSSI nch_mac L=30N W=220N M=1
MN5 QAB AWT2 NET46 VSSI nch_mac L=30N W=300N M=1
MN6 NET46 NET085 VSSI VSSI nch_mac L=30N W=300N M=1
MM33 NET0144 SEL_AB NET0205 VSSI nch_mac L=30N W=220N M=1
MM0 NET130 GBL VSSI VSSI nch_mac L=30N W=300N M=3
MN21 QBB_T QB_T NET130 VSSI nch_mac L=30N W=300N M=3
MM25 QB_T QBB_T Z3 VSSI nch_mac L=30N W=330N M=3
MM53 QAB QB_T NET0142 VDDI pch_mac L=30N W=440N M=1
MM50 NET0210 AWT2 VDDI VDDI pch_mac L=30N W=300N M=1
MM47 NET0192 SEL_B NET0210 VDDI pch_mac L=30N W=300N M=1
MM46 NET0194 SEL_BB VDDI VDDI pch_mac L=30N W=0.88U M=3
MM45 QBB QBBB NET0192 VDDI pch_mac L=30N W=300N M=1
MM38 NET069 AWT1B QBB VDDI pch_mac L=30N W=300N M=2
MM48 NET0206 AWT2 VDDI VDDI pch_mac L=30N W=300N M=1
MM54 QBB QB_T NET0194 VDDI pch_mac L=30N W=0.5U M=3
MM39 NET069 NET0173 VDDI VDDI pch_mac L=30N W=300N M=2
MM44 QBB QB_T NET0194 VDDI pch_mac L=30N W=440N M=1
MP4 QBB_T QB_T VDDI VDDI pch_mac L=30N W=880N M=1
MM35 NET0141 SEL_A NET0206 VDDI pch_mac L=30N W=300N M=1
MM30 QAB QB_T NET0142 VDDI pch_mac L=30N W=0.5U M=3
MP10 NET48 AWT1B QAB VDDI pch_mac L=30N W=300N M=2
MP11 NET48 NET085 VDDI VDDI pch_mac L=30N W=300N M=2
MP7 VDDI DLRSB GBLB VDDI pch_mac L=30N W=1U M=6
MP0 GBLB GBL VDDI VDDI pch_mac L=30N W=320N M=1
MM29 NET0142 SEL_AB VDDI VDDI pch_mac L=30N W=0.88U M=3
MP6 VDDI GBLB GBL VDDI pch_mac L=30N W=320N M=1
MM34 QAB QABB NET0141 VDDI pch_mac L=30N W=300N M=1
MP8 GBL DLRSB VDDI VDDI pch_mac L=30N W=1U M=6
MM28 QB_T QBB_T VDDI VDDI pch_mac L=30N W=880N M=1
MM27 QB_T GBLB VDDI VDDI pch_mac L=30N W=880N M=1
MP15 QBB_T GBL VDDI VDDI pch_mac L=30N W=0.88U M=2
XI210 AWT QLATCH_BB VSSI VSSI VDDI VDDI SEL_B SDBM200W80_NOR_BULK FN1=1 WN1=0.3U 
+ LN1=0.03U FN2=1 WN2=0.3U LN2=0.03U FP2=1 WP2=0.5U LP2=0.03U MULTI=1 FP1=2 
+ WP1=0.5U LP1=0.03U
XI174 AWT QLATCH_AB VSSI VSSI VDDI VDDI SEL_A SDBM200W80_NOR_BULK FN1=1 WN1=0.3U 
+ LN1=0.03U FN2=1 WN2=0.3U LN2=0.03U FP2=1 WP2=0.5U LP2=0.03U MULTI=1 FP1=2 
+ WP1=0.5U LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    LPLCH_DE_DATA
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_LPLCH_DE_DATA CKC CKT IN Q QB VDDI VSSI
*.PININFO CKC:I CKT:I IN:I Q:O QB:O VDDI:B VSSI:B
MM3 NET037 CKT VSSI VSSI nch_mac L=30N W=150N M=1
MM2 QB Q NET037 VSSI nch_mac L=30N W=150N M=1
MM11 QB IN NET38 VSSI nch_mac L=30N W=210N M=1
MM8 NET38 CKC VSSI VSSI nch_mac L=30N W=210N M=1
MM1 QB Q NET036 VDDI pch_mac L=30N W=150N M=1
MM0 NET036 CKC VDDI VDDI pch_mac L=30N W=150N M=1
MM9 NET39 CKT VDDI VDDI pch_mac L=30N W=320N M=1
MM10 QB IN NET39 VDDI pch_mac L=30N W=320N M=1
XI1 QB VSSI VSSI VDDI VDDI Q SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 FP=1 
+ WP=0.32U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    PHASE_SEL_DATA
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_PHASE_SEL_DATA PHASE1 PHASE2 SEL SELB SELOUT VDDI VSSI
*.PININFO PHASE1:I PHASE2:I SEL:I SELB:I SELOUT:B VDDI:B VSSI:B
MM11 SELOUT SEL NET08 VSSI nch_mac L=30N W=320N M=1
MM8 NET08 PHASE2 VSSI VSSI nch_mac L=30N W=320N M=1
MM5 SELOUT SELB NET015 VSSI nch_mac L=30N W=320N M=1
MM4 NET015 PHASE1 VSSI VSSI nch_mac L=30N W=320N M=1
MM10 SELOUT SELB NET038 VDDI pch_mac L=30N W=540N M=1
MM9 NET038 PHASE2 VDDI VDDI pch_mac L=30N W=540N M=1
MM7 NET039 PHASE1 VDDI VDDI pch_mac L=30N W=540N M=1
MM6 SELOUT SEL NET039 VDDI pch_mac L=30N W=540N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DIN_MUX_V1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DIN_MUX_V1 AWTDA AWTDB BWEBA BWEBABX BWEBB DA DABX DB DCLK PHASESEL 
+ VDDI VSSI
*.PININFO BWEBA:I BWEBB:I DA:I DB:I DCLK:I PHASESEL:I AWTDA:O AWTDB:O 
*.PININFO BWEBABX:O DABX:O VDDI:B VSSI:B
XI17 CKC CKT BWEBBX2 BWEBBXT BWEBBXC VDDI VSSI SDBM200W80_LPLCH_DE_DATA
XDB_LATCH CKC CKT DBX2 DBXT DBXC VDDI VSSI SDBM200W80_LPLCH_DE_DATA
XI28 SELB VSSI VSSI VDDI VDDI SEL SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI27 PHASESEL VSSI VSSI VDDI VDDI SELB SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.32U LP=0.03U
XI16 BWEBBX1B VSSI VSSI VDDI VDDI BWEBBX2 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI15 BWEBB VSSI VSSI VDDI VDDI BWEBBX1B SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI12 BWEBAX1B VSSI VSSI VDDI VDDI BWEBAX2 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI11 BWEBA VSSI VSSI VDDI VDDI BWEBAX1B SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI10 DBX1B VSSI VSSI VDDI VDDI DBX2 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 
+ FP=1 WP=0.21U LP=0.03U
XI9 DB VSSI VSSI VDDI VDDI DBX1B SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 
+ FP=1 WP=0.21U LP=0.03U
XI8 DAX1B VSSI VSSI VDDI VDDI DAX2 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 
+ FP=1 WP=0.21U LP=0.03U
XI7 DA VSSI VSSI VDDI VDDI DAX1B SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 
+ FP=1 WP=0.21U LP=0.03U
XI4 CKC VSSI VSSI VDDI VDDI CKT SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 FP=1 
+ WP=0.32U LP=0.03U
XI3 DCLK VSSI VSSI VDDI VDDI CKC SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XBWEB_MUX BWEBAX2 BWEBBXT SEL SELB BWEBABX VDDI VSSI SDBM200W80_PHASE_SEL_DATA
XD_MUX DAX2 DBXT SEL SELB DABX VDDI VSSI SDBM200W80_PHASE_SEL_DATA
MM4 ZB20 BWEBBX1B VSSI VSSI nch_mac L=30N W=150N M=1
MM5 ZB20 DBX2 VSSI VSSI nch_mac L=30N W=150N M=1
MM6 AWTDB BWEBBX2 ZB20 VSSI nch_mac L=30N W=150N M=1
MM7 AWTDB DBX1B ZB20 VSSI nch_mac L=30N W=150N M=1
MN6 AWTDA DAX1B ZA20 VSSI nch_mac L=30N W=150N M=1
MN13 ZA20 DAX2 VSSI VSSI nch_mac L=30N W=150N M=1
MN4 ZA20 BWEBAX1B VSSI VSSI nch_mac L=30N W=150N M=1
MN5 AWTDA BWEBAX2 ZA20 VSSI nch_mac L=30N W=150N M=1
MM8 AWTDB DBX1B NET21 VDDI pch_mac L=30N W=210N M=1
MM9 AWTDB DBX2 NET25 VDDI pch_mac L=30N W=210N M=1
MM10 NET25 BWEBBX1B VDDI VDDI pch_mac L=30N W=210N M=1
MM11 NET21 BWEBBX2 VDDI VDDI pch_mac L=30N W=210N M=1
MP5 AWTDA DAX2 NET17 VDDI pch_mac L=30N W=210N M=1
MP4 NET17 BWEBAX1B VDDI VDDI pch_mac L=30N W=210N M=1
MP3 NET13 BWEBAX2 VDDI VDDI pch_mac L=30N W=210N M=1
MP2 AWTDA DAX1B NET13 VDDI pch_mac L=30N W=210N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    IO_WOBIST_DP
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_IO_WOBIST_DP AWT BWEBA BWEBB CKD DA DB DCLK DCLKA GBL GBLB GW GWB 
+ PHASESEL QA QB QLATCH_AB QLATCH_BB RSC_TRK_W VDDI VSSI WLP_SAEB
*.PININFO AWT:I BWEBA:I BWEBB:I CKD:I DA:I DB:I DCLK:I DCLKA:I PHASESEL:I 
*.PININFO QLATCH_AB:I QLATCH_BB:I WLP_SAEB:I GW:O GWB:O QA:O QB:O GBL:B GBLB:B 
*.PININFO RSC_TRK_W:B VDDI:B VSSI:B
XDIN BWEBABX CKD DABX DCLKA GW GWB VDDI VSSI SDBM200W80_DIN_WOBIST_DP_V2
XDOUT AWT AWTDA AWTDB GBL GBLB QA QB QLATCH_AB QLATCH_BB VDDI VSSI WLP_SAEB 
+ SDBM200W80_DOUT_DP_V1
XDIN_MUX AWTDA AWTDB BWEBA BWEBABX BWEBB DA DABX DB DCLK PHASESEL VDDI VSSI 
+ SDBM200W80_DIN_MUX_V1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    PRECHARGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_PRECHARGE BL BLB BLEQB VDDI
*.PININFO BLEQB:I BL:B BLB:B VDDI:B
MP0_MIXV_SLH VDDI BLEQB BL VDDI pch_mac L=30N W=0.44U M=3
MP5_MIXV_SLH BL BLEQB BLB VDDI pch_mac L=30N W=440N M=1
MP17_MIXV_SLH BLB BLEQB VDDI VDDI pch_mac L=30N W=0.44U M=3
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    YPASS_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_YPASS_M4 BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] BLEQ 
+ BLEQB DL DLB VDDI VSSI WC WT Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
*.PININFO BLEQ:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I Y[6]:I Y[7]:I 
*.PININFO BLEQB:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B 
*.PININFO BLB[3]:B DL:B DLB:B VDDI:B VSSI:B WC:B WT:B
XI1 BLEQ VSSI VSSI VDDI VDDI NET37 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.21U LP=0.03U
XI[0] Y[0] VSSI VSSI VDDI VDDI YB[0] SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
XI[1] Y[1] VSSI VSSI VDDI VDDI YB[1] SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
XI[2] Y[2] VSSI VSSI VDDI VDDI YB[2] SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
XI[3] Y[3] VSSI VSSI VDDI VDDI YB[3] SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
MM2[0] BLB[0] BL[0] VDDI VDDI pch_mac L=30N W=120N M=1
MM2[1] BLB[1] BL[1] VDDI VDDI pch_mac L=30N W=120N M=1
MM2[2] BLB[2] BL[2] VDDI VDDI pch_mac L=30N W=120N M=1
MM2[3] BLB[3] BL[3] VDDI VDDI pch_mac L=30N W=120N M=1
MM3[0] BL[0] BLB[0] VDDI VDDI pch_mac L=30N W=120N M=1
MM3[1] BL[1] BLB[1] VDDI VDDI pch_mac L=30N W=120N M=1
MM3[2] BL[2] BLB[2] VDDI VDDI pch_mac L=30N W=120N M=1
MM3[3] BL[3] BLB[3] VDDI VDDI pch_mac L=30N W=120N M=1
MP0 VDDI BLEQB DL VDDI pch_mac L=30N W=150N M=1
MP10[0] DLB YB[0] BLB[0] VDDI pch_mac L=30N W=370N M=1
MP10[1] DLB YB[1] BLB[1] VDDI pch_mac L=30N W=370N M=1
MP10[2] DLB YB[2] BLB[2] VDDI pch_mac L=30N W=370N M=1
MP10[3] DLB YB[3] BLB[3] VDDI pch_mac L=30N W=370N M=1
MP2 DLB BLEQB VDDI VDDI pch_mac L=30N W=150N M=1
MM1 BLEQB NET37 VDDI VDDI pch_mac L=30N W=1.12U M=1
MP1[0] DL YB[0] BL[0] VDDI pch_mac L=30N W=370N M=1
MP1[1] DL YB[1] BL[1] VDDI pch_mac L=30N W=370N M=1
MP1[2] DL YB[2] BL[2] VDDI pch_mac L=30N W=370N M=1
MP1[3] DL YB[3] BL[3] VDDI pch_mac L=30N W=370N M=1
MM0 BLEQB NET37 VSSI VSSI nch_mac L=30N W=245N M=2
MN31_MIXV_SLS[0] BL[0] Y[4] WT VSSI nch_mac L=30N W=820N M=1
MN31_MIXV_SLS[1] BL[1] Y[5] WT VSSI nch_mac L=30N W=820N M=1
MN31_MIXV_SLS[2] BL[2] Y[6] WT VSSI nch_mac L=30N W=820N M=1
MN31_MIXV_SLS[3] BL[3] Y[7] WT VSSI nch_mac L=30N W=820N M=1
MN30_MIXV_SLS[0] BLB[0] Y[4] WC VSSI nch_mac L=30N W=820N M=1
MN30_MIXV_SLS[1] BLB[1] Y[5] WC VSSI nch_mac L=30N W=820N M=1
MN30_MIXV_SLS[2] BLB[2] Y[6] WC VSSI nch_mac L=30N W=820N M=1
MN30_MIXV_SLS[3] BLB[3] Y[7] WC VSSI nch_mac L=30N W=820N M=1
XPRECHARGE[0] BL[0] BLB[0] BLEQB VDDI SDBM200W80_PRECHARGE
XPRECHARGE[1] BL[1] BLB[1] BLEQB VDDI SDBM200W80_PRECHARGE
XPRECHARGE[2] BL[2] BLB[2] BLEQB VDDI SDBM200W80_PRECHARGE
XPRECHARGE[3] BL[3] BLB[3] BLEQB VDDI SDBM200W80_PRECHARGE
.ENDS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    NAND_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_NAND_BULK A B G GB P PB Y
*.PININFO A:I B:I G:I GB:I P:I PB:I Y:O
M1 Y A P PB pch_mac L=LP1 W=WP1 M=MULTI*FP1
M4 Y B P PB pch_mac L=LP2 W=WP2 M=MULTI*FP2
M6 Y B NET9 GB nch_mac L=LN2 W=WN2 M=MULTI*FN2
M8 NET9 A G GB nch_mac L=LN1 W=WN1 M=MULTI*FN1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    SA_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_SA_M4 DLB_DN DLB_UP DL_DN DL_UP GBL GBLB PGB_DN PGB_UP PREB SAE VDDI 
+ VSSI
*.PININFO PGB_DN:I PGB_UP:I PREB:I SAE:I DLB_DN:B DLB_UP:B DL_DN:B DL_UP:B 
*.PININFO GBL:B GBLB:B VDDI:B VSSI:B
MN0 DL_IN DLB_IN NS VSSI nch_mac L=90N W=0.5U M=4
MN2 NS SAE VSSI VSSI nch_mac L=30N W=0.5U M=4
MN1 DLB_IN DL_IN NS VSSI nch_mac L=90N W=0.5U M=4
MN11 GBL SO VSSI VSSI nch_mac L=35.0N W=0.67U M=6
MN12 GBLB SOB VSSI VSSI nch_mac L=35.0N W=0.67U M=6
MP2 DL_IN DLB_IN VDDI VDDI pch_mac L=30N W=500N M=1
MP10 DL_IN PREB VDDI VDDI pch_mac L=30N W=500N M=1
MP6 DL_UP PGB_UP DL_IN VDDI pch_mac L=30N W=500N M=1
MP14 DLB_IN PGB_DN DLB_DN VDDI pch_mac L=30N W=500N M=1
MP7 DLB_IN PGB_UP DLB_UP VDDI pch_mac L=30N W=500N M=1
MP13 DL_DN PGB_DN DL_IN VDDI pch_mac L=30N W=500N M=1
MP3 DLB_IN DL_IN VDDI VDDI pch_mac L=30N W=500N M=1
MP8 DL_IN PREB DLB_IN VDDI pch_mac L=30N W=500N M=2
MP11 DLB_IN PREB VDDI VDDI pch_mac L=30N W=500N M=1
XINV1 DLB_IN VSSI VSSI VDDI VDDI SOB SDBM200W80_INV_BULK FN=1 WN=0.2U LN=0.03U MULTI=1 
+ FP=3 WP=0.22U LP=0.03U
XINV0 DL_IN VSSI VSSI VDDI VDDI SO SDBM200W80_INV_BULK FN=1 WN=0.2U LN=0.03U MULTI=1 
+ FP=3 WP=0.22U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    NAND3_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_NAND3_BULK A B C G GB P PB Y
*.PININFO A:I B:I C:I G:I GB:I P:I PB:I Y:O
M1 Y A P PB pch_mac L=LP1 W=WP1 M=MULTI*FP1
M3 Y B P PB pch_mac L=LP2 W=WP2 M=MULTI*FP2
M7 Y C P PB pch_mac L=LP3 W=WP3 M=MULTI*FP3
M9 Y C NET17 GB nch_mac L=LN3 W=WN3 M=MULTI*FN3
M11 NET17 B NET14 GB nch_mac L=LN2 W=WN2 M=MULTI*FN2
M13 NET14 A G GB nch_mac L=LN1 W=WN1 M=MULTI*FN1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    IO_RWBLK_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_IO_RWBLK_M4 BLEQB_DN BLEQB_UP BLEQ_DN BLEQ_UP DLB_DN DLB_UP DL_DN 
+ DL_UP GBL GBLB GW GWB PREBG SAEB VDDI VSSI WC WT
*.PININFO BLEQB_DN:I BLEQB_UP:I BLEQ_DN:I BLEQ_UP:I GW:I GWB:I PREBG:I SAEB:I 
*.PININFO WC:O WT:O DLB_DN:B DLB_UP:B DL_DN:B DL_UP:B GBL:B GBLB:B VDDI:B 
*.PININFO VSSI:B
MP25 WT GWB VDDI VDDI pch_mac L=30N W=0.21U M=5
MP27 WC GW VDDI VDDI pch_mac L=30N W=0.21U M=5
MN0 WC GW VSSI VSSI nch_mac L=30N W=0.49U M=7
MN13 WT GWB VSSI VSSI nch_mac L=30N W=0.49U M=7
XI222 SAEC PREBGB VSSI VSSI VDDI VDDI PREB SDBM200W80_NAND_BULK FN1=1 WN1=0.25U 
+ LN1=0.03U FN2=1 WN2=0.25U LN2=0.03U FP2=1 WP2=0.32U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.32U LP1=0.03U
XSA DLB_DN DLB_UP DL_DN DL_UP GBL GBLB PGB_DN PGB_UP PREB SAE VDDI VSSI SDBM200W80_SA_M4
XI38 BLEQB_UP VSSI VSSI VDDI VDDI PGB_UP SDBM200W80_INV_BULK FN=1 WN=0.24U LN=0.03U 
+ MULTI=1 FP=1 WP=0.36U LP=0.03U
XI37 BLEQB_DN VSSI VSSI VDDI VDDI PGB_DN SDBM200W80_INV_BULK FN=1 WN=0.24U LN=0.03U 
+ MULTI=1 FP=1 WP=0.36U LP=0.03U
XI54 PREBG VSSI VSSI VDDI VDDI PREBGB SDBM200W80_INV_BULK FN=1 WN=0.25U LN=0.03U 
+ MULTI=1 FP=1 WP=0.32U LP=0.03U
XI248 SAEC VSSI VSSI VDDI VDDI SAE SDBM200W80_INV_BULK FN=1 WN=0.16U LN=0.03U MULTI=1 
+ FP=1 WP=0.33U LP=0.03U
XI235 GBLB GBL SAEB VSSI VSSI VDDI VDDI SAEC SDBM200W80_NAND3_BULK FN1=1 WN1=0.29U 
+ LN1=0.03U FN2=1 WN2=0.29U LN2=0.03U FN3=1 WN3=0.29U LN3=0.03U FP3=1 
+ WP3=0.16U LP3=0.03U FP2=1 WP2=0.16U LP2=0.03U MULTI=1 FP1=1 WP1=0.16U 
+ LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    YPASS_M4_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_YPASS_M4_D BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] BLEQ 
+ BLEQB DL DLB VDDI VSSI WC WT Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
*.PININFO BLEQ:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I Y[6]:I Y[7]:I 
*.PININFO BLEQB:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B 
*.PININFO BLB[3]:B DL:B DLB:B VDDI:B VSSI:B WC:B WT:B
XI1 BLEQ VSSI VSSI VDDI VDDI NET37 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.21U LP=0.03U
XI[0] Y[0] VSSI VSSI VDDI VDDI YB[0] SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
XI[1] Y[1] VSSI VSSI VDDI VDDI YB[1] SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
XI[2] Y[2] VSSI VSSI VDDI VDDI YB[2] SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
XI[3] Y[3] VSSI VSSI VDDI VDDI YB[3] SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
MM2[0] BLB[0] BL[0] VDDI VDDI pch_mac L=30N W=120N M=1
MM2[1] BLB[1] BL[1] VDDI VDDI pch_mac L=30N W=120N M=1
MM2[2] BLB[2] BL[2] VDDI VDDI pch_mac L=30N W=120N M=1
MM2[3] BLB[3] BL[3] VDDI VDDI pch_mac L=30N W=120N M=1
MM3[0] BL[0] BLB[0] VDDI VDDI pch_mac L=30N W=120N M=1
MM3[1] BL[1] BLB[1] VDDI VDDI pch_mac L=30N W=120N M=1
MM3[2] BL[2] BLB[2] VDDI VDDI pch_mac L=30N W=120N M=1
MM3[3] BL[3] BLB[3] VDDI VDDI pch_mac L=30N W=120N M=1
MP0 VDDI BLEQB DL VDDI pch_mac L=30N W=150N M=1
MP10[0] DLB YB[0] BLB[0] VDDI pch_mac L=30N W=370N M=1
MP10[1] DLB YB[1] BLB[1] VDDI pch_mac L=30N W=370N M=1
MP10[2] DLB YB[2] BLB[2] VDDI pch_mac L=30N W=370N M=1
MP10[3] DLB YB[3] BLB[3] VDDI pch_mac L=30N W=370N M=1
MP2 DLB BLEQB VDDI VDDI pch_mac L=30N W=150N M=1
MM1 BLEQB NET37 VDDI VDDI pch_mac L=30N W=1.12U M=1
MP1[0] DL YB[0] BL[0] VDDI pch_mac L=30N W=370N M=1
MP1[1] DL YB[1] BL[1] VDDI pch_mac L=30N W=370N M=1
MP1[2] DL YB[2] BL[2] VDDI pch_mac L=30N W=370N M=1
MP1[3] DL YB[3] BL[3] VDDI pch_mac L=30N W=370N M=1
MM0 BLEQB NET37 VSSI VSSI nch_mac L=30N W=490N M=1
MN31_MIXV_SLS[0] BL[0] Y[4] WT VSSI nch_mac L=30N W=820N M=1
MN31_MIXV_SLS[1] BL[1] Y[5] WT VSSI nch_mac L=30N W=820N M=1
MN31_MIXV_SLS[2] BL[2] Y[6] WT VSSI nch_mac L=30N W=820N M=1
MN31_MIXV_SLS[3] BL[3] Y[7] WT VSSI nch_mac L=30N W=820N M=1
MN30_MIXV_SLS[0] BLB[0] Y[4] WC VSSI nch_mac L=30N W=820N M=1
MN30_MIXV_SLS[1] BLB[1] Y[5] WC VSSI nch_mac L=30N W=820N M=1
MN30_MIXV_SLS[2] BLB[2] Y[6] WC VSSI nch_mac L=30N W=820N M=1
MN30_MIXV_SLS[3] BLB[3] Y[7] WC VSSI nch_mac L=30N W=820N M=1
XPRECHARGE[0] BL[0] BLB[0] BLEQB VDDI SDBM200W80_PRECHARGE
XPRECHARGE[1] BL[1] BLB[1] BLEQB VDDI SDBM200W80_PRECHARGE
XPRECHARGE[2] BL[2] BLB[2] BLEQB VDDI SDBM200W80_PRECHARGE
XPRECHARGE[3] BL[3] BLB[3] BLEQB VDDI SDBM200W80_PRECHARGE
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    LIO_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_LIO_M4 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_UP[0] BLB_UP[1] 
+ BLB_UP[2] BLB_UP[3] BLEQ_DN BLEQ_UP BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] 
+ BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] GBL GBLB GW GWB PREBG SAEB VDDI VSSI 
+ Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] 
+ Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I PREBG:I SAEB:I Y_DN[0]:I Y_DN[1]:I 
*.PININFO Y_DN[2]:I Y_DN[3]:I Y_DN[4]:I Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I 
*.PININFO Y_UP[0]:I Y_UP[1]:I Y_UP[2]:I Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I 
*.PININFO Y_UP[6]:I Y_UP[7]:I BLB_DN[0]:B BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B 
*.PININFO BLB_UP[0]:B BLB_UP[1]:B BLB_UP[2]:B BLB_UP[3]:B BL_DN[0]:B 
*.PININFO BL_DN[1]:B BL_DN[2]:B BL_DN[3]:B BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B 
*.PININFO BL_UP[3]:B GBL:B GBLB:B VDDI:B VSSI:B
XYPASS_U BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BLB_UP[0] BLB_UP[1] BLB_UP[2] 
+ BLB_UP[3] BLEQ_UP BLEQB_UP_0 DL_UP DLB_UP VDDI VSSI WC WT Y_UP[0] Y_UP[1] 
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_YPASS_M4
XIO_RWBLK BLEQB_DN_0 BLEQB_UP_0 BLEQ_DN BLEQ_UP DLB_DN DLB_UP DL_DN DL_UP GBL 
+ GBLB GW GWB PREBG SAEB VDDI VSSI WC WT SDBM200W80_IO_RWBLK_M4
XYPASS_D BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BLB_DN[0] BLB_DN[1] BLB_DN[2] 
+ BLB_DN[3] BLEQ_DN BLEQB_DN_0 DL_DN DLB_DN VDDI VSSI WC WT Y_DN[0] Y_DN[1] 
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] SDBM200W80_YPASS_M4_D
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    XDRV_WLP_M
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_XDRV_WLP_M BLEQ BLEQB BS BSB DEC_X2[0] DEC_X2[1] VDDI VSSI WLPY[0] 
+ WLPY[1]
*.PININFO BS:I DEC_X2[0]:I DEC_X2[1]:I BLEQ:O BLEQB:O BSB:O WLPY[0]:O 
*.PININFO WLPY[1]:O VDDI:B VSSI:B
XI534 MWL2[0] VSSI VSSI VDDI VDDI WLPY[0] SDBM200W80_INV_BULK FN=3 WN=1.5U LN=0.03U 
+ MULTI=1 FP=6 WP=1.5U LP=0.03U
XI532 NET022 VSSI VSSI VDDI VDDI WLPY[1] SDBM200W80_INV_BULK FN=3 WN=1.5U LN=0.03U 
+ MULTI=1 FP=6 WP=1.5U LP=0.03U
XI557 BSB VSSI VSSI VDDI VDDI BLEQ SDBM200W80_INV_BULK FN=6 WN=0.7U LN=0.03U MULTI=1 
+ FP=6 WP=0.9U LP=0.03U
XI595 BSB VSSI VSSI VDDI VDDI BLEQB SDBM200W80_INV_BULK FN=2 WN=0.9U LN=0.03U MULTI=1 
+ FP=2 WP=1.2U LP=0.03U
XI551 BS VSSI VSSI VDDI VDDI BSB SDBM200W80_INV_BULK FN=1 WN=0.9U LN=0.03U MULTI=1 FP=1 
+ WP=1.2U LP=0.03U
MM9 NET022 BS VDDI VDDI pch_mac L=30N W=0.7U M=3
MM20 MWL2[0] BS VDDI VDDI pch_mac L=30N W=0.7U M=3
MM12 MWL2[0] DEC_X2[0] VDDI VDDI pch_mac L=30N W=350N M=2
MM10 NET022 DEC_X2[1] VDDI VDDI pch_mac L=30N W=350N M=2
MM0 SHARE BS VSSI VSSI nch_mac L=30N W=1U M=6
MM32 NET022 DEC_X2[1] SHARE VSSI nch_mac L=30N W=0.7U M=5
MM28 MWL2[0] DEC_X2[0] SHARE VSSI nch_mac L=30N W=0.7U M=5
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    XDRV_Y4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_XDRV_Y4 VDDI VSSI WLPY YIN[0] YIN[1] YIN[2] YIN[3] YOUT[0] YOUT[1] 
+ YOUT[2] YOUT[3]
*.PININFO WLPY:I YIN[0]:I YIN[1]:I YIN[2]:I YIN[3]:I YOUT[0]:O YOUT[1]:O 
*.PININFO YOUT[2]:O YOUT[3]:O VDDI:B VSSI:B
MM34 YOUT[3] MWL2[3] VSSI VSSI nch_mac L=30N W=0.73U M=8
MM31 MWL2[3] YIN[3] SHARE VSSI nch_mac L=30N W=0.72U M=4
MM28 MWL2[2] YIN[2] SHARE VSSI nch_mac L=30N W=0.72U M=4
MM23 YOUT[1] MWL2[1] VSSI VSSI nch_mac L=30N W=0.73U M=8
MM26 YOUT[2] MWL2[2] VSSI VSSI nch_mac L=30N W=0.73U M=8
MM2 MWL2[0] YIN[0] SHARE VSSI nch_mac L=30N W=0.72U M=4
MM5 YOUT[0] MWL2[0] VSSI VSSI nch_mac L=30N W=0.73U M=8
MN21 SHARE WLPY VSSI VSSI nch_mac L=30N W=0.8U M=8
MM21 MWL2[1] YIN[1] SHARE VSSI nch_mac L=30N W=0.72U M=4
MM1 MWL2[0] YIN[0] VDDI VDDI pch_mac L=30N W=0.68U M=3
MM24 YOUT[1] MWL2[1] VDDI VDDI pch_mac L=30N W=0.8U M=14
MM3 MWL2[0] WLPY VDDI VDDI pch_mac L=30N W=0.68U M=3
MM25 YOUT[2] MWL2[2] VDDI VDDI pch_mac L=30N W=0.8U M=14
MP31 SHARE WLPY VDDI VDDI pch_mac L=30N W=150N M=2
MM4 YOUT[0] MWL2[0] VDDI VDDI pch_mac L=30N W=0.8U M=14
MM32 MWL2[3] YIN[3] VDDI VDDI pch_mac L=30N W=0.68U M=3
MM30 MWL2[2] WLPY VDDI VDDI pch_mac L=30N W=0.68U M=3
MM20 MWL2[1] WLPY VDDI VDDI pch_mac L=30N W=0.68U M=3
MM33 MWL2[3] WLPY VDDI VDDI pch_mac L=30N W=0.68U M=3
MM35 YOUT[3] MWL2[3] VDDI VDDI pch_mac L=30N W=0.8U M=14
MM27 MWL2[2] YIN[2] VDDI VDDI pch_mac L=30N W=0.68U M=3
MM22 MWL2[1] YIN[1] VDDI VDDI pch_mac L=30N W=0.68U M=3
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    XDRV_READ
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_XDRV_READ BS SAEB VDDI VSSI WLP_SAE
*.PININFO BS:I WLP_SAE:I SAEB:O VDDI:B VSSI:B
XNAND0_MIXV_SLH BS WLP_SAE VSSI VSSI VDDI VDDI BS_WLPSAEB SDBM200W80_NAND_BULK FN1=2 
+ WN1=0.75U LN1=0.03U FN2=2 WN2=0.75U LN2=0.03U FP2=2 WP2=0.45U LP2=0.03U 
+ MULTI=1 FP1=2 WP1=0.45U LP1=0.03U
XI426_MIXV_SLH BS_WLPSAEB VSSI VSSI VDDI VDDI SAEB SDBM200W80_INV_BULK FN=4 WN=0.9U 
+ LN=0.03U MULTI=1 FP=7 WP=1U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    LCTRL_M
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_LCTRL_M BLEQB_DN BLEQB_UP BSB_DN BSB_UP DEC_X3_DN DEC_X3_UP DEC_Y[0] 
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] 
+ DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] 
+ DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] 
+ DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] PREBG SAEB VDDI VSSI WLP_SAE
*.PININFO BLEQB_DN:I BLEQB_UP:I BSB_DN:I BSB_UP:I DEC_X3_DN:I DEC_X3_UP:I 
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I WLP_SAE:I DEC_Y_DN[0]:O DEC_Y_DN[1]:O 
*.PININFO DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O DEC_Y_DN[5]:O 
*.PININFO DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O DEC_Y_UP[1]:O 
*.PININFO DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O DEC_Y_UP[5]:O 
*.PININFO DEC_Y_UP[6]:O DEC_Y_UP[7]:O PREBG:O SAEB:O VDDI:B VSSI:B
XNOR0_MIXV_SLH DEC_X3_UP DEC_X3_DN VSSI VSSI VDDI VDDI BS0 SDBM200W80_NOR_BULK FN1=1 
+ WN1=0.4U LN1=0.03U FN2=1 WN2=0.4U LN2=0.03U FP2=1 WP2=0.7U LP2=0.03U MULTI=1 
+ FP1=1 WP1=0.7U LP1=0.03U
XXDRV_Y4_D[0] VDDI VSSI BLEQB_DN DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] SDBM200W80_XDRV_Y4
XXDRV_Y4_D[1] VDDI VSSI BLEQB_DN DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] SDBM200W80_XDRV_Y4
XXDRV_Y4_U[0] VDDI VSSI BLEQB_UP DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] SDBM200W80_XDRV_Y4
XXDRV_Y4_U[1] VDDI VSSI BLEQB_UP DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] SDBM200W80_XDRV_Y4
XI251 BSB_UP BSB_DN VSSI VSSI VDDI VDDI NET0105 SDBM200W80_NAND_BULK FN1=1 WN1=0.87U 
+ LN1=0.03U FN2=1 WN2=0.87U LN2=0.03U FP2=1 WP2=0.54U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.54U LP1=0.03U
XNAND0_MIXV_SLH BS0 BS5 VSSI VSSI VDDI VDDI NET28 SDBM200W80_NAND_BULK FN1=1 WN1=0.4U 
+ LN1=0.03U FN2=1 WN2=0.4U LN2=0.03U FP2=1 WP2=0.75U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.75U LP1=0.03U
XXDRV_READ BSD SAEB VDDI VSSI WLP_SAE SDBM200W80_XDRV_READ
XINV4_MIXV_SLH BS4 VSSI VSSI VDDI VDDI BS4B SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV5_MIXV_SLH BS4B VSSI VSSI VDDI VDDI BS5 SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XI253 NET0105 VSSI VSSI VDDI VDDI NET0102 SDBM200W80_INV_BULK FN=2 WN=0.65U LN=0.03U 
+ MULTI=1 FP=2 WP=0.87U LP=0.03U
XI254 NET0102 VSSI VSSI VDDI VDDI PREBG SDBM200W80_INV_BULK FN=6 WN=0.87U LN=0.03U 
+ MULTI=1 FP=8 WP=0.87U LP=0.03U
XI249 NET28 VSSI VSSI VDDI VDDI NET93 SDBM200W80_INV_BULK FN=1 WN=0.16U LN=0.03U 
+ MULTI=1 FP=1 WP=0.16U LP=0.03U
XI250 NET93 VSSI VSSI VDDI VDDI BSD SDBM200W80_INV_BULK FN=1 WN=0.16U LN=0.03U MULTI=1 
+ FP=1 WP=0.16U LP=0.03U
XINV0_MIXV_SLH BS0 VSSI VSSI VDDI VDDI BS1B SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV3_MIXV_SLH BS3B VSSI VSSI VDDI VDDI BS4 SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV2_MIXV_SLH BS2 VSSI VSSI VDDI VDDI BS3B SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV1_MIXV_SLH BS1B VSSI VSSI VDDI VDDI BS2 SDBM200W80_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    LCTRL_M_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_LCTRL_M_M4 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] 
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] 
+ DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] 
+ DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] PREBG SAEB VDDI 
+ VSSI WLPY_DN[0] WLPY_DN[1] WLPY_UP[0] WLPY_UP[1] WLP_SAE WLP_SAE_TK
*.PININFO BLEQ_DN:O BLEQ_UP:O DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O 
*.PININFO DEC_Y_DN[3]:O DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O 
*.PININFO DEC_Y_DN[7]:O DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O 
*.PININFO DEC_Y_UP[3]:O DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O 
*.PININFO DEC_Y_UP[7]:O PREBG:O SAEB:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_UP[0]:O 
*.PININFO WLPY_UP[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X3[0]:B 
*.PININFO DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B 
*.PININFO DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B 
*.PININFO DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B VDDI:B VSSI:B WLP_SAE:B 
*.PININFO WLP_SAE_TK:B
XXDRV_WLP_DN BLEQ_DN BLEQB_DN DEC_X3[0] BSB_DN DEC_X2[0] DEC_X2[1] VDDI VSSI 
+ WLPY_DN[0] WLPY_DN[1] SDBM200W80_XDRV_WLP_M
XXDRV_WLP_UP BLEQ_UP BLEQB_UP DEC_X3[1] BSB_UP DEC_X2[0] DEC_X2[1] VDDI VSSI 
+ WLPY_UP[0] WLPY_UP[1] SDBM200W80_XDRV_WLP_M
XLCTRL BLEQB_DN BLEQB_UP BSB_DN BSB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] 
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] 
+ DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] 
+ DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] 
+ DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] PREBG SAEB VDDI VSSI WLP_SAE SDBM200W80_LCTRL_M
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    XDRV_STRAP_LCNT
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_XDRV_STRAP_LCNT VDDI VSSI WLPY WLPYB
*.PININFO WLPY:I VDDI:B VSSI:B WLPYB:B
MN1 WLPYB WLPY VSSI VSSI nch_mac L=30N W=2U M=4
MP0 WLPYB WLPY VDDI VDDI pch_mac L=30N W=1.8U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    XDRV_LA512_SHA
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_XDRV_LA512_SHA DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] SH_NPD VDDI VSSI WLOUT[0] WLOUT[1] WLPY WLPYB WLP_SAE 
+ WLP_SAE_TK
*.PININFO WLPY:I WLPYB:I WLP_SAE:I WLOUT[0]:O WLOUT[1]:O DEC_X0[0]:B 
*.PININFO DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B 
*.PININFO DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B 
*.PININFO DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B 
*.PININFO DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B DEC_X3[0]:B 
*.PININFO DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B 
*.PININFO DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B 
*.PININFO DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B SH_NPD:B VDDI:B VSSI:B 
*.PININFO WLP_SAE_TK:B
MP20_MIXV_SLH WLOUT[0] MWL2 VDDI VDDI pch_mac L=35.0N W=1.15U M=6
MP7 MWL0 DEC_X1[0] VDDI VDDI pch_mac L=35.0N W=150N M=1
MP14 MWL0A DEC_X0[1] VDDI VDDI pch_mac L=35.0N W=150N M=1
MM1_MIXV_SLH WLOUT[1] MWL2A VDDI VDDI pch_mac L=35.0N W=1.15U M=6
MM3 VDDI WLPY MWL2A VDDI pch_mac L=35.0N W=0.64U M=2
MM8 MWL2 MWL1 VDDI VDDI pch_mac L=35.0N W=0.5U M=2
MM5 MWL2A MWL1A VDDI VDDI pch_mac L=35.0N W=0.5U M=2
MP19 VDDI WLPY MWL2 VDDI pch_mac L=35.0N W=0.64U M=2
MP13 MWL0A DEC_X1[0] VDDI VDDI pch_mac L=35.0N W=150N M=1
MP6 MWL0 DEC_X0[0] VDDI VDDI pch_mac L=35.0N W=150N M=1
MN7 MWL0A DEC_X0[1] SH_NPD VSSI nch_mac L=35.0N W=150N M=1
MN0 MWL2 MWL1 WLPYB VSSI nch_mac L=35.0N W=0.9U M=2
MP9 MWL0 DEC_X0[0] SH_NPD VSSI nch_mac L=35.0N W=150N M=1
MM2_MIXV_SLH WLOUT[1] MWL2A VSSI VSSI nch_mac L=35.0N W=1U M=4
MM4 MWL2A MWL1A WLPYB VSSI nch_mac L=35.0N W=0.9U M=2
MN6_MIXV_SLH WLOUT[0] MWL2 VSSI VSSI nch_mac L=35.0N W=1U M=4
XI426 MWL0A VSSI VSSI VDDI VDDI MWL1A SDBM200W80_INV_BULK FN=1 WN=0.39U LN=0.03U 
+ MULTI=1 FP=1 WP=0.565U LP=0.03U
XI425 MWL0 VSSI VSSI VDDI VDDI MWL1 SDBM200W80_INV_BULK FN=1 WN=0.39U LN=0.03U MULTI=1 
+ FP=1 WP=0.565U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    XDRV_LA512_SHA_NMOS
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_XDRV_LA512_SHA_NMOS DEC_X1 SH_NPD VSSI
*.PININFO DEC_X1:B SH_NPD:B VSSI:B
MN5 SH_NPD DEC_X1 VSSI VSSI nch_mac L=35.0N W=320N M=2
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TKBL_TRKPRE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TKBL_TRKPRE TRKBL TRKWL VDDI VSSI ZH ZL
*.PININFO TRKWL:I ZH:O ZL:O TRKBL:B VDDI:B VSSI:B
MM7 ZH NET_021 VDDI VDDI pch_mac L=30N W=0.98U M=3
MM8 NET_039 NET_039 VDDI VDDI pch_mac L=30N W=210N M=2
MP0_MIXV_SLH TRKBL TRKWL VDDI VDDI pch_mac L=30N W=1.2U M=3
MM4 NET_039 NET_021 VDDI VDDI pch_mac L=30N W=210N M=2
MM01 ZL NET_039 VSSI VSSI nch_mac L=30N W=1.09U M=3
MM2 NET_021 NET_021 VSSI VSSI nch_mac L=30N W=210N M=2
MM3 NET_021 NET_039 VSSI VSSI nch_mac L=30N W=210N M=2
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TKBL_EDGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TKBL_EDGE BLB_EDGE BL_EDGE G_FLOAT VDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I BLB_EDGE:B BL_EDGE:B G_FLOAT:B VDDI:B VSSI:B TIEH:B
MPCHPU1 BLB TIEH VDDI VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDI BLB TIEH VDDI pchpu_sr L=35N W=40N M=1
MNCHPD1 BLB TIEH VSSI VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 G_FLOAT BLB TIEH VSSI nchpd_sr L=35N W=95N M=1
MNCHPG1 BLB WL BL_EDGE VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 BLB_EDGE WL TIEH VSSI nchpg_sr L=35N W=65N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TKBL_BCELL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TKBL_BCELL BLB BL_TK G_FLOAT VDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I BLB:B BL_TK:B G_FLOAT:B VDDI:B VSSI:B TIEH:B
MPCHPU1 TIEH BL_TK_IN VDDI VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDI TIEH BL_TK_IN VDDI pchpu_sr L=35N W=40N M=1
MNCHPD1 TIEH BL_TK_IN G_FLOAT VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 VSSI TIEH BL_TK_IN VSSI nchpd_sr L=35N W=95N M=1
MNCHPG1 TIEH WL BLB VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 BL_TK WL_TK BL_TK_IN VSSI nchpg_sr L=35N W=65N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TRKNOR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TRKNOR BLB BLB_EDGE BL_EDGE BL_TK G_FLOAT VDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I TIEH:I BLB:B BLB_EDGE:B BL_EDGE:B BL_TK:B G_FLOAT:B 
*.PININFO VDDI:B VSSI:B
XTKBL_BCELL_RIGHT BLB_EDGE BL_EDGE G_FLOAT VDDI VSSI WL WL_TK TIEH SDBM200W80_TKBL_EDGE
XTKBL_BCELL BLB BL_TK G_FLOAT VDDI VSSI WL WL_TK TIEH SDBM200W80_TKBL_BCELL
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TRKNORX2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TRKNORX2 BL_TK VDDI VSSI WL[0] WL[1] WL_TK FLOAT1 FLOAT2 FLOAT3 FLOAT4 
+ FLOAT5 TIEH
*.PININFO WL[0]:I WL[1]:I WL_TK:I TIEH:I BL_TK:B VDDI:B VSSI:B FLOAT1:B 
*.PININFO FLOAT2:B FLOAT3:B FLOAT4:B FLOAT5:B
XTRKNOR_1 FLOAT2 FLOAT4 FLOAT1 BL_TK G_FLOAT VDDI VSSI WL[1] WL_TK TIEH 
+ SDBM200W80_TRKNOR
XTRKNOR_0 FLOAT3 FLOAT5 FLOAT1 BL_TK G_FLOAT VDDI VSSI WL[0] WL_TK TIEH 
+ SDBM200W80_TRKNOR
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    MCB_TKWL_ISO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_MCB_TKWL_ISO BL BLB VDDI VSSI WLL WLR
*.PININFO BL:B BLB:B VDDI:B VSSI:B WLL:B WLR:B
MNCHPG1 BLB WLR VSSI VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 NET060 WLL BL VSSI nchpg_sr L=35N W=65N M=1
MNCHPD1 VSSI NET060 VSSI VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 VSSI VSSI NET060 VSSI nchpd_sr L=35N W=95N M=1
MPCHPU1 VSSI NET060 P_FLOAT VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDI VSSI NET060 VDDI pchpu_sr L=35N W=40N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    MCB_TKWL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_MCB_TKWL BL BLB VDDI VSSI WL
*.PININFO BL:B BLB:B VDDI:B VSSI:B WL:B
MPCHPU1 VSSI BL_IN P_FLOAT VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDI VSSI BL_IN VDDI pchpu_sr L=35N W=40N M=1
MNCHPD1 VSSI BL_IN VSSI VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 VSSI VSSI BL_IN VSSI nchpd_sr L=35N W=95N M=1
MNCHPG1 BLB WL VSSI VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 BL_IN WL BL VSSI nchpg_sr L=35N W=65N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TKWL_2X2_ISO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TKWL_2X2_ISO VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] WL_TK_R[1]
*.PININFO WL_TK_L[0]:I WL_TK_L[1]:I WL_TK_R[0]:I WL_TK_R[1]:I VDDI:B VSSI:B
XI24 NET030 NET284 VDDI VSSI WL_TK_R[0] SDBM200W80_MCB_TKWL
XTKWL_MCB_1 NET281 NET284 VDDI VSSI WL_TK_R[1] SDBM200W80_MCB_TKWL
XI25 NET294 NET278 VDDI VSSI WL_TK_R[0] WL_TK_L[0] SDBM200W80_MCB_TKWL_ISO
XI22 NET279 NET278 VDDI VSSI WL_TK_R[1] WL_TK_L[1] SDBM200W80_MCB_TKWL_ISO
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TKWL_2X2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TKWL_2X2 VDDI VSSI WL_DUM WL_TK
*.PININFO VDDI:B VSSI:B WL_DUM:B WL_TK:B
XTKWL_MCB_1 FLOAT_BL_R_T FLOAT_BLB_R VDDI VSSI WL_TK SDBM200W80_MCB_TKWL
XTKWL_MCB_0 FLOAT_BL_L_T FLOAT_BLB_L VDDI VSSI WL_TK SDBM200W80_MCB_TKWL
XTKDUM_MCB_1 FLOAT_BL_R_B FLOAT_BLB_R VDDI VSSI WL_DUM SDBM200W80_MCB_TKWL
XTKDUM_MCB_0 FLOAT_BL_L_B FLOAT_BLB_L VDDI VSSI WL_DUM SDBM200W80_MCB_TKWL
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    MCB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_MCB BL BLB VDDI VSSI WL
*.PININFO BL:B BLB:B VDDI:B VSSI:B WL:B
MPCHPU1 BLB_IN BL_IN VDDI VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDI BLB_IN BL_IN VDDI pchpu_sr L=35N W=40N M=1
MNCHPD1 BLB_IN BL_IN VSSI VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 VSSI BLB_IN BL_IN VSSI nchpd_sr L=35N W=95N M=1
MNCHPG1 BLB WL BLB_IN VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 BL_IN WL BL VSSI nchpg_sr L=35N W=65N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    MCB_2X4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_MCB_2X4 BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB 
+ GW GWB VDDI VSSI WL[0] WL[1]
*.PININFO BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B 
*.PININFO GBL:B GBLB:B GW:B GWB:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XMCB_0[0] BL[0] BLB[0] VDDI VSSI WL[0] SDBM200W80_MCB
XMCB_0[1] BL[1] BLB[1] VDDI VSSI WL[0] SDBM200W80_MCB
XMCB_0[2] BL[2] BLB[2] VDDI VSSI WL[0] SDBM200W80_MCB
XMCB_0[3] BL[3] BLB[3] VDDI VSSI WL[0] SDBM200W80_MCB
XMCB_1[0] BL[0] BLB[0] VDDI VSSI WL[1] SDBM200W80_MCB
XMCB_1[1] BL[1] BLB[1] VDDI VSSI WL[1] SDBM200W80_MCB
XMCB_1[2] BL[2] BLB[2] VDDI VSSI WL[1] SDBM200W80_MCB
XMCB_1[3] BL[3] BLB[3] VDDI VSSI WL[1] SDBM200W80_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DIO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DIO A VSSI
*.PININFO A:B VSSI:B
DDIO VSSI A ndio AREA=0.02E-12 M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TOP_EDGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TOP_EDGE VDDI VSSI WLP_SAE WLP_SAE_TK
*.PININFO VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XI58 NET023 VSSI VSSI VDDI VDDI WLP_SAE_TK SDBM200W80_INV_BULK FN=9 WN=0.8U LN=0.03U 
+ MULTI=1 FP=16 WP=0.675U LP=0.03U
XI55 WLP_SAE VSSI VSSI VDDI VDDI NET023 SDBM200W80_INV_BULK FN=3 WN=0.9U LN=0.03U 
+ MULTI=1 FP=3 WP=1.2U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CLK_BUF_DP_V2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CLK_BUF_DP_V2 CKC CKPB1_L CKPB_EN CKT VDDI VSSI WCLK_L WCLK_R
*.PININFO CKPB1_L:I CKPB_EN:I CKC:O CKT:O WCLK_L:O WCLK_R:O VDDI:B VSSI:B
XI1 CKPB1_L CKPB_EN VSSI VSSI VDDI VDDI NET42 SDBM200W80_NAND_BULK FN1=2 WN1=0.98U 
+ LN1=0.03U FN2=2 WN2=0.98U LN2=0.03U FP2=2 WP2=0.76U LP2=0.03U MULTI=1 FP1=2 
+ WP1=0.76U LP1=0.03U
XI2 NET050 VSSI VSSI VDDI VDDI NET51 SDBM200W80_INV_BULK FN=2 WN=0.76U LN=0.03U MULTI=1 
+ FP=2 WP=0.98U LP=0.03U
XI28 CKC VSSI VSSI VDDI VDDI CKT SDBM200W80_INV_BULK FN=3 WN=0.76U LN=0.03U MULTI=1 
+ FP=3 WP=0.98U LP=0.03U
XI9 NET51 VSSI VSSI VDDI VDDI WCLK_R SDBM200W80_INV_BULK FN=5 WN=0.76U LN=0.03U MULTI=1 
+ FP=5 WP=0.98U LP=0.03U
XI10 NET51 VSSI VSSI VDDI VDDI WCLK_L SDBM200W80_INV_BULK FN=5 WN=0.76U LN=0.03U 
+ MULTI=1 FP=5 WP=0.98U LP=0.03U
XI3 NET42 VSSI VSSI VDDI VDDI CKC SDBM200W80_INV_BULK FN=3 WN=0.76U LN=0.03U MULTI=1 
+ FP=3 WP=0.98U LP=0.03U
XI5 NET051 VSSI VSSI VDDI VDDI NET050 SDBM200W80_INV_BULK FN=1 WN=0.76U LN=0.03U 
+ MULTI=1 FP=1 WP=0.98U LP=0.03U
XI4 NET42 VSSI VSSI VDDI VDDI NET051 SDBM200W80_INV_BULK FN=1 WN=0.76U LN=0.03U MULTI=1 
+ FP=1 WP=0.98U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    N_AORBANDC
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_N_AORBANDC A B C OUT VDDI VSSI
*.PININFO A:I B:I C:I OUT:O VDDI:B VSSI:B
MM8 OUT C NET13 VSSI nch_mac L=30N W=540N M=1
MM7 NET13 A VSSI VSSI nch_mac L=30N W=540N M=1
MM6 NET13 B VSSI VSSI nch_mac L=30N W=540N M=1
MM11 NET27 A VDDI VDDI pch_mac L=30N W=650N M=1
MM10 OUT B NET27 VDDI pch_mac L=30N W=650N M=1
MM9 OUT C VDDI VDDI pch_mac L=30N W=430N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CKP_GEN_DOUBLE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CKP_GEN_DOUBLE CE CKPB CKP_RSTB CLK CLK2 VDDI VSSI
*.PININFO CE:I CKP_RSTB:I CLK:I CLK2:I CKPB:O VDDI:B VSSI:B
MM12 NET41 CKPBB NET81 VSSI nch_mac L=30N W=540N M=1
MM10 NET81 CKP_RSTB VSSI VSSI nch_mac L=30N W=540N M=1
MM9 CKPB CLK_ENB2 NET41 VSSI nch_mac L=30N W=540N M=1
MM8 CKPB CLKB2 NET41 VSSI nch_mac L=30N W=540N M=1
MM0 NET83 CLK_EN VSSI VSSI nch_mac L=30N W=0.98U M=3
MM18 CKPB CLK NET83 VSSI nch_mac L=30N W=0.98U M=2
MM7 CKPB CLKB2 NET82 VDDI pch_mac L=30N W=0.98U M=2
MM6 NET82 CLK_ENB2 VDDI VDDI pch_mac L=30N W=0.98U M=3
MM3 CKPB CLK_EN NET74 VDDI pch_mac L=30N W=540N M=1
MM2 NET74 CKPBB VDDI VDDI pch_mac L=30N W=540N M=1
MM1 NET74 CKP_RSTB VDDI VDDI pch_mac L=30N W=540N M=1
MM15 CKPB CLK NET74 VDDI pch_mac L=30N W=540N M=1
XI20 CLK_EN2 VSSI VSSI VDDI VDDI CLK_ENB2 SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U 
+ MULTI=1 FP=1 WP=0.43U LP=0.03U
XI22 NET84 VSSI VSSI VDDI VDDI CLK_EN2 SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U 
+ MULTI=1 FP=1 WP=0.43U LP=0.03U
XI21 CE VSSI VSSI VDDI VDDI NET56 SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U MULTI=1 
+ FP=1 WP=0.54U LP=0.03U
XI8 CKPBB VSSI VSSI VDDI VDDI NET53 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI7 CLK VSSI VSSI VDDI VDDI NET85 SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U MULTI=1 
+ FP=1 WP=0.54U LP=0.03U
XI2 CKPB VSSI VSSI VDDI VDDI CKPBB SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI17 CLK2 VSSI VSSI VDDI VDDI CLKB2 SDBM200W80_INV_BULK FN=1 WN=0.54U LN=0.03U MULTI=1 
+ FP=1 WP=0.87U LP=0.03U
XI3 CLK_ENB NET56 VSSI VSSI VDDI VDDI CLK_EN SDBM200W80_NOR_BULK FN1=1 WN1=0.32U 
+ LN1=0.03U FN2=1 WN2=0.32U LN2=0.03U FP2=1 WP2=0.54U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.54U LP1=0.03U
XI18 CLK_EN2 CLKB2 CKPBB NET84 VDDI VSSI SDBM200W80_N_AORBANDC
XI10 CLK_EN NET85 NET53 CLK_ENB VDDI VSSI SDBM200W80_N_AORBANDC
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    RESETD_TSEL_WT_NEW
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_RESETD_TSEL_WT_NEW CKPB VDDI VSSI OUT WV[0] WV[1]
*.PININFO CKPB:I WV[0]:I WV[1]:I OUT:O VDDI:B VSSI:B
XI91 NET36 WV[1] VSSI VSSI VDDI VDDI NET46 SDBM200W80_NAND_BULK FN1=1 WN1=0.32U 
+ LN1=0.03U FN2=1 WN2=0.32U LN2=0.03U FP2=1 WP2=0.21U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.21U LP1=0.03U
XI90 NET12 NET46 VSSI VSSI VDDI VDDI OUT SDBM200W80_NAND_BULK FN1=1 WN1=0.32U LN1=0.03U 
+ FN2=1 WN2=0.32U LN2=0.03U FP2=1 WP2=0.21U LP2=0.03U MULTI=1 FP1=1 WP1=0.21U 
+ LP1=0.03U
MM11 NET60 NET33 VDDI VDDI pch_mac L=30N W=150N M=1
MM10 NET36 NET33 NET60 VDDI pch_mac L=30N W=150N M=1
MM1 NET12 CKPB NET64 VDDI pch_mac L=30N W=320N M=1
MM0 NET12 WV[0] VDDI VDDI pch_mac L=30N W=210N M=1
MM31 NET64 Z4 VDDI VDDI pch_mac L=30N W=320N M=1
MM15 Z4 NET46 NET58 VDDI pch_mac L=30N W=150N M=1
MM5 NET33 CKPB NET63 VDDI pch_mac L=30N W=150N M=1
MM14 NET58 NET46 VDDI VDDI pch_mac L=30N W=150N M=1
MM4 NET63 CKPB VDDI VDDI pch_mac L=30N W=150N M=1
MM9 NET36 NET33 NET61 VSSI nch_mac L=30N W=150N M=1
MM3 NET12 Z4 NET15 VSSI nch_mac L=30N W=320N M=1
MM2 NET12 CKPB NET15 VSSI nch_mac L=30N W=320N M=1
MM22 NET15 WV[0] VSSI VSSI nch_mac L=30N W=320N M=1
MM8 NET61 NET33 VSSI VSSI nch_mac L=30N W=150N M=1
MM13 NET59 NET46 VSSI VSSI nch_mac L=30N W=150N M=1
MM7 NET62 CKPB VSSI VSSI nch_mac L=30N W=150N M=1
MM6 NET33 CKPB NET62 VSSI nch_mac L=30N W=150N M=1
MM12 Z4 NET46 NET59 VSSI nch_mac L=30N W=150N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    PTSEL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_PTSEL CKP2LOW_TSEL[0] CKP2LOW_TSEL[1] IN OUT VDDI VSSI
*.PININFO CKP2LOW_TSEL[0]:I CKP2LOW_TSEL[1]:I IN:I OUT:B VDDI:B VSSI:B
XI7 IN VSSI VSSI VDDI VDDI NET21 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U MULTI=1 
+ FP=1 WP=0.65U LP=0.03U
XTSEL_DWL_LOW NET21 VDDI VSSI NET045 CKP2LOW_TSEL[0] CKP2LOW_TSEL[1] 
+ SDBM200W80_RESETD_TSEL_WT_NEW
XI1 NET045 NET21 VSSI VSSI VDDI VDDI OUT SDBM200W80_NOR_BULK FN1=4 WN1=0.65U LN1=0.03U 
+ FN2=4 WN2=0.65U LN2=0.03U FP2=4 WP2=1.2U LP2=0.03U MULTI=1 FP1=4 WP1=1.2U 
+ LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CKPB2_GEN_V2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CKPB2_GEN_V2 AT CE CKPB CLK RSC VDDI VSSI
*.PININFO AT:I CE:I CLK:I RSC:I CKPB:O VDDI:B VSSI:B
XI7 CLK VSSI VSSI VDDI VDDI NET57 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI2 CKPB VSSI VSSI VDDI VDDI NET51 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI8 NET51 VSSI VSSI VDDI VDDI NET31 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI9 NET57 CLK_EN NET31 NET56 VDDI VSSI SDBM200W80_N_AORBANDC
XI3 NET56 AT VSSI VSSI VDDI VDDI CLK_EN SDBM200W80_NOR_BULK FN1=1 WN1=0.54U LN1=0.03U 
+ FN2=1 WN2=0.54U LN2=0.03U FP2=1 WP2=0.98U LP2=0.03U MULTI=1 FP1=1 WP1=0.98U 
+ LP1=0.03U
MM18 CKPB CLK NET59 VSSI nch_mac L=30N W=0.98U M=5
MM0 NET59 CLK_EN VSSI VSSI nch_mac L=30N W=0.98U M=6
MM4 CKPB NET51 NET58 VSSI nch_mac L=30N W=980N M=1
MM5 NET58 RSC VSSI VSSI nch_mac L=30N W=980N M=1
MM14 CKPB NET51 NET45 VDDI pch_mac L=30N W=980N M=1
MM15 CKPB RSC NET45 VDDI pch_mac L=30N W=0.98U M=5
MM16 NET45 CLK_EN VDDI VDDI pch_mac L=30N W=0.98U M=7
MM1 NET45 CLK VDDI VDDI pch_mac L=30N W=980N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CKPB1_GEN_V1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CKPB1_GEN_V1 AT CE CKPB CLK RSC VDDI VSSI
*.PININFO AT:I CE:I CLK:I RSC:I CKPB:O VDDI:B VSSI:B
MM5 NET74 RSC VSSI VSSI nch_mac L=30N W=980N M=1
MM4 CKPB NET68 NET74 VSSI nch_mac L=30N W=980N M=1
MM0 NET76 CLK_EN VSSI VSSI nch_mac L=30N W=0.98U M=6
MM18 CKPB CLK NET76 VSSI nch_mac L=30N W=0.98U M=5
MM14 CKPB NET68 NET66 VDDI pch_mac L=30N W=980N M=1
MM16 NET66 CLK_EN VDDI VDDI pch_mac L=30N W=0.98U M=7
MM1 NET66 CLK VDDI VDDI pch_mac L=30N W=980N M=1
MM15 CKPB RSC NET66 VDDI pch_mac L=30N W=0.98U M=5
XI8 NET68 VSSI VSSI VDDI VDDI NET073 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI7 CLK VSSI VSSI VDDI VDDI NET069 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI2 CKPB VSSI VSSI VDDI VDDI NET68 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI3 NET034 CE VSSI VSSI VDDI VDDI CLK_EN SDBM200W80_NOR_BULK FN1=1 WN1=0.65U LN1=0.03U 
+ FN2=1 WN2=0.65U LN2=0.03U FP2=1 WP2=0.98U LP2=0.03U MULTI=1 FP1=1 WP1=0.98U 
+ LP1=0.03U
XI9 NET069 CLK_EN NET073 NET034 VDDI VSSI SDBM200W80_N_AORBANDC
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CKG_GEN_V7
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CKG_GEN_V7 CEAI CEBAI CEBBI CEBI CKP1 CKP2 CKP2SEL[0] CKP2SEL[1] CKPB1 
+ CKPB1_TRK CKPB2 CKPB_EN CKP_EN CKP_RSTB CKTA CLK TIE_H VDDI VSSI
*.PININFO CEAI:I CEBAI:I CEBBI:I CEBI:I CKP2SEL[0]:I CKP2SEL[1]:I CKP_RSTB:I 
*.PININFO CKTA:I CLK:I TIE_H:I CKP1:O CKP2:O CKPB1:O CKPB1_TRK:O CKPB2:O 
*.PININFO CKPB_EN:O CKP_EN:O VDDI:B VSSI:B
XI41 NET66 CKPB2 NET0142 VSSI VSSI VDDI VDDI CKP_EN_RSTB SDBM200W80_NAND3_BULK FN1=1 
+ WN1=0.76U LN1=0.03U FN2=1 WN2=0.76U LN2=0.03U FN3=1 WN3=0.76U LN3=0.03U 
+ FP3=1 WP3=0.32U LP3=0.03U FP2=1 WP2=0.32U LP2=0.03U MULTI=1 FP1=1 WP1=0.32U 
+ LP1=0.03U
XI6 CEAI CEBI VSSI VSSI VDDI VDDI CE SDBM200W80_NOR_BULK FN1=1 WN1=0.43U LN1=0.03U 
+ FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.98U LP2=0.03U MULTI=1 FP1=1 WP1=0.98U 
+ LP1=0.03U
XI19 NET0157 CKP_RST3 VSSI VSSI VDDI VDDI NET66 SDBM200W80_NOR_BULK FN1=1 WN1=0.32U 
+ LN1=0.03U FN2=1 WN2=0.32U LN2=0.03U FP2=1 WP2=0.65U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.65U LP1=0.03U
XI14 CKP_RSTB2_TRK CKP_RSTB4_TRK VSSI VSSI VDDI VDDI CKP_RST3 SDBM200W80_NAND_BULK 
+ FN1=1 WN1=0.65U LN1=0.03U FN2=1 WN2=0.65U LN2=0.03U FP2=1 WP2=0.32U 
+ LP2=0.03U MULTI=1 FP1=1 WP1=0.32U LP1=0.03U
XI13 CKP_RSTB CKPB1_TRK VSSI VSSI VDDI VDDI NET0157 SDBM200W80_NAND_BULK FN1=1 
+ WN1=0.43U LN1=0.03U FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.32U LP2=0.03U 
+ MULTI=1 FP1=1 WP1=0.32U LP1=0.03U
XSELECT_GEN CEBI CKPB_EN CKP_EN_RSTB CKPB1_TRK_5D CKPB2 VDDI VSSI 
+ SDBM200W80_CKP_GEN_DOUBLE
XI12 CKPB1_TRK VSSI VSSI VDDI VDDI NET0145 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI144 CKPB1 VSSI VSSI VDDI VDDI CKP1 SDBM200W80_INV_BULK FN=3 WN=0.65U LN=0.03U MULTI=1 
+ FP=3 WP=0.87U LP=0.03U
XI129 CKPB_EN VSSI VSSI VDDI VDDI CKP_EN SDBM200W80_INV_BULK FN=5 WN=0.76U LN=0.03U 
+ MULTI=1 FP=5 WP=0.98U LP=0.03U
XI77 NET0134 VSSI VSSI VDDI VDDI CKP_RSTB3 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI79 CKPB2 VSSI VSSI VDDI VDDI CKP2 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U MULTI=1 
+ FP=1 WP=0.65U LP=0.03U
XI3 NET0117 VSSI VSSI VDDI VDDI CKPB1_TRK_5D SDBM200W80_INV_BULK FN=1 WN=0.54U LN=0.03U 
+ MULTI=1 FP=1 WP=0.76U LP=0.03U
XI24 NET0168 VSSI VSSI VDDI VDDI NET0142 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI2 NET0156 VSSI VSSI VDDI VDDI NET0117 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI18 CKP2 VSSI VSSI VDDI VDDI NET0167 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI20 NET0167 VSSI VSSI VDDI VDDI NET0168 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
MM25 NET0227 NET0145 VSSI VSSI nch_mac L=30N W=160N M=1
MM9 NET0151 NET0145 NET0227 VSSI nch_mac L=30N W=160N M=1
MM33 NET0225 NET0151 VSSI VSSI nch_mac L=30N W=160N M=1
MM34 NET0156 NET0151 NET0225 VSSI nch_mac L=30N W=160N M=1
MM40 NET0134 NET0129 NET0160 VSSI nch_mac L=30N W=150N M=1
MM41 NET0160 NET0129 VSSI VSSI nch_mac L=30N W=150N M=1
MM32 NET0129 NET0130 NET0146 VSSI nch_mac L=30N W=150N M=1
MM37 NET0146 NET0130 VSSI VSSI nch_mac L=30N W=150N M=1
MM49 NET0153 CKP_RSTB2_TRK VSSI VSSI nch_mac L=30N W=150N M=1
MM29 NET0149 CKP_RSTB4_TRK VSSI VSSI nch_mac L=30N W=150N M=1
MM28 NET0130 CKP_RSTB4_TRK NET0149 VSSI nch_mac L=30N W=150N M=1
MM46 CKP_RSTB4_TRK NET0153 VSSI VSSI nch_mac L=30N W=150N M=1
MM26 NET0151 NET0145 VDDI VDDI pch_mac L=30N W=160N M=1
MM36 NET0156 NET0151 VDDI VDDI pch_mac L=30N W=160N M=1
MM42 NET0144 NET0129 VDDI VDDI pch_mac L=30N W=150N M=1
MM43 NET0134 NET0129 NET0144 VDDI pch_mac L=30N W=150N M=1
MM39 NET0129 NET0130 NET0147 VDDI pch_mac L=30N W=150N M=1
MM38 NET0147 NET0130 VDDI VDDI pch_mac L=30N W=150N M=1
MM31 NET0130 CKP_RSTB4_TRK NET0148 VDDI pch_mac L=30N W=150N M=1
MM30 NET0148 CKP_RSTB4_TRK VDDI VDDI pch_mac L=30N W=150N M=1
MM52 CKP_RSTB4_TRK NET0153 VDDI VDDI pch_mac L=30N W=150N M=1
MM48 NET0153 CKP_RSTB2_TRK VDDI VDDI pch_mac L=30N W=150N M=1
XI10 CKP2SEL[0] CKP2SEL[1] CKP_RSTB CKP_RSTB2_TRK VDDI VSSI SDBM200W80_PTSEL
XCKPB2_GEN CKPB_EN CEBBI CKPB2 CKP_RSTB2_TRK CKP_RSTB VDDI VSSI SDBM200W80_CKPB2_GEN_V2
XCKPB1_GEN_TRK TIE_H CE CKPB1_TRK CLK CKP_RSTB VDDI VSSI SDBM200W80_CKPB1_GEN_V1
XCKPB1_GEN TIE_H CEBAI CKPB1 CLK CKP_RSTB VDDI VSSI SDBM200W80_CKPB1_GEN_V1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    Q_LATCH_CLK_1007
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_Q_LATCH_CLK_1007 CEBAF CKPB1 CKPB2 CKP_RSTB CKTA CKTA2 IOSAE QCLKBA_L 
+ QCLKBA_R QCLKBB_L QCLKBB_R VDDI VSSI
*.PININFO CEBAF:I CKPB1:I CKPB2:I CKP_RSTB:I IOSAE:I CKTA:O CKTA2:O QCLKBA_L:O 
*.PININFO QCLKBA_R:O QCLKBB_L:O QCLKBB_R:O VDDI:B VSSI:B
XI12 NET0132 IOSAE VSSI VSSI VDDI VDDI NET0168 SDBM200W80_NAND_BULK FN1=2 WN1=0.98U 
+ LN1=0.03U FN2=2 WN2=0.98U LN2=0.03U FP2=2 WP2=0.76U LP2=0.03U MULTI=1 FP1=2 
+ WP1=0.76U LP1=0.03U
XI5 NET0113 IOSAE VSSI VSSI VDDI VDDI NET049 SDBM200W80_NAND_BULK FN1=2 WN1=0.98U 
+ LN1=0.03U FN2=2 WN2=0.98U LN2=0.03U FP2=2 WP2=0.76U LP2=0.03U MULTI=1 FP1=2 
+ WP1=0.76U LP1=0.03U
MM3 NET0119 IOSAE NET0171 VSSI nch_mac L=30N W=120N M=1
MM1 NET0171 NET0132 VSSI VSSI nch_mac L=30N W=120N M=1
MM19 NET0112 CKTA2 NET0128 VSSI nch_mac L=30N W=210N M=1
MM20 NET0112 IOSAE NET0126 VSSI nch_mac L=30N W=120N M=1
MM49 NET0128 IOSAEB VSSI VSSI nch_mac L=30N W=210N M=1
MM21 NET0126 NET0113 VSSI VSSI nch_mac L=30N W=120N M=1
MM2 NET0119 CKTB2 NET0172 VSSI nch_mac L=30N W=210N M=1
MM0 NET0172 IOSAEB VSSI VSSI nch_mac L=30N W=210N M=1
XI35 NET0206 VSSI VSSI VDDI VDDI NET0205 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI34 NET0207 VSSI VSSI VDDI VDDI NET0204 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI33 CKTA VSSI VSSI VDDI VDDI NET0206 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI14 NET0159 VSSI VSSI VDDI VDDI QCLKBB_L SDBM200W80_INV_BULK FN=5 WN=0.76U LN=0.03U 
+ MULTI=1 FP=5 WP=0.98U LP=0.03U
XI13 NET0159 VSSI VSSI VDDI VDDI QCLKBB_R SDBM200W80_INV_BULK FN=5 WN=0.76U LN=0.03U 
+ MULTI=1 FP=5 WP=0.98U LP=0.03U
XI11 NET0119 VSSI VSSI VDDI VDDI NET0132 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U 
+ MULTI=1 FP=1 WP=0.65U LP=0.03U
XI10 NET0168 VSSI VSSI VDDI VDDI NET0159 SDBM200W80_INV_BULK FN=2 WN=0.76U LN=0.03U 
+ MULTI=1 FP=2 WP=0.98U LP=0.03U
XI20 NET0179 VSSI VSSI VDDI VDDI NET0177 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI24 NET0190 VSSI VSSI VDDI VDDI NET0189 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI23 NET0189 VSSI VSSI VDDI VDDI CKTB2 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.32U LP=0.03U
XI22 CKCB VSSI VSSI VDDI VDDI NET0190 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI3 NET0112 VSSI VSSI VDDI VDDI NET0113 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U 
+ MULTI=1 FP=1 WP=0.65U LP=0.03U
XI32 CKTB VSSI VSSI VDDI VDDI NET0207 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI15 IOSAE VSSI VSSI VDDI VDDI IOSAEB SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U 
+ MULTI=1 FP=1 WP=0.43U LP=0.03U
XI27 NET0204 VSSI VSSI VDDI VDDI CKCB SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI21 NET0177 VSSI VSSI VDDI VDDI CKTA2 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.32U LP=0.03U
XI30 NET30 VSSI VSSI VDDI VDDI QCLKBA_R SDBM200W80_INV_BULK FN=5 WN=0.76U LN=0.03U 
+ MULTI=1 FP=5 WP=0.98U LP=0.03U
XI29 NET30 VSSI VSSI VDDI VDDI QCLKBA_L SDBM200W80_INV_BULK FN=5 WN=0.76U LN=0.03U 
+ MULTI=1 FP=5 WP=0.98U LP=0.03U
XI26 CKPB2 VSSI VSSI VDDI VDDI CKTB SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI18 CKPB1 VSSI VSSI VDDI VDDI CKTA SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XI25 NET0205 VSSI VSSI VDDI VDDI CKCA SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
XI7 NET049 VSSI VSSI VDDI VDDI NET30 SDBM200W80_INV_BULK FN=2 WN=0.76U LN=0.03U MULTI=1 
+ FP=2 WP=0.98U LP=0.03U
XI19 CKCA VSSI VSSI VDDI VDDI NET0179 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U 
+ MULTI=1 FP=1 WP=0.15U LP=0.03U
MM7 NET0169 NET0132 VDDI VDDI pch_mac L=30N W=120N M=1
MM6 NET0170 IOSAE VDDI VDDI pch_mac L=30N W=320N M=1
MM5 NET0119 IOSAEB NET0169 VDDI pch_mac L=30N W=120N M=1
MM4 NET0119 CKTB2 NET0170 VDDI pch_mac L=30N W=320N M=1
MM26 NET0112 IOSAEB NET0125 VDDI pch_mac L=30N W=120N M=1
MM29 NET0112 CKTA2 NET0127 VDDI pch_mac L=30N W=320N M=1
MM50 NET0127 IOSAE VDDI VDDI pch_mac L=30N W=320N M=1
MM51 NET0125 NET0113 VDDI VDDI pch_mac L=30N W=120N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    LPLCH_CEB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_LPLCH_CEB CKC CKT IN Q QB VDDI VSSI
*.PININFO CKC:I CKT:I IN:I Q:O QB:O VDDI:B VSSI:B
MM3 NET037 CKT VSSI VSSI nch_mac L=30N W=120N M=1
MM2 NET023 Q NET037 VSSI nch_mac L=30N W=120N M=1
MM11 NET023 IN NET38 VSSI nch_mac L=30N W=430N M=1
MM8 NET38 CKC VSSI VSSI nch_mac L=30N W=430N M=1
MM1 NET023 Q NET036 VDDI pch_mac L=30N W=120N M=1
MM0 NET036 CKC VDDI VDDI pch_mac L=30N W=120N M=1
MM9 NET39 CKT VDDI VDDI pch_mac L=30N W=540N M=1
MM10 NET023 IN NET39 VDDI pch_mac L=30N W=540N M=1
XI2 Q VSSI VSSI VDDI VDDI QB SDBM200W80_INV_BULK FN=1 WN=0.65U LN=0.03U MULTI=1 FP=1 
+ WP=0.87U LP=0.03U
XI1 NET023 VSSI VSSI VDDI VDDI Q SDBM200W80_INV_BULK FN=1 WN=0.65U LN=0.03U MULTI=1 
+ FP=1 WP=0.87U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    PHASE_SEL_ADD_V1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_PHASE_SEL_ADD_V1 PHASE1 PHASE2 SEL1B SEL2 SELOUT VDDI VSSI
*.PININFO PHASE1:I PHASE2:I SEL1B:I SEL2:I SELOUT:B VDDI:B VSSI:B
MM11 SELOUT SEL2 NET08 VSSI nch_mac L=30N W=430N M=1
MM8 NET08 PHASE2 VSSI VSSI nch_mac L=30N W=430N M=1
MM5 SELOUT SEL1B NET015 VSSI nch_mac L=30N W=540N M=1
MM4 NET015 PHASE1 VSSI VSSI nch_mac L=30N W=540N M=1
MM10 SELOUT SEL1B NET038 VDDI pch_mac L=30N W=540N M=1
MM9 NET038 PHASE2 VDDI VDDI pch_mac L=30N W=540N M=1
MM7 NET039 PHASE1 VDDI VDDI pch_mac L=30N W=760N M=1
MM6 SELOUT SEL2 NET039 VDDI pch_mac L=30N W=760N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    LPLCH_DE_ADD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_LPLCH_DE_ADD CKC CKT IN Q QB VDDI VSSI
*.PININFO CKC:I CKT:I IN:I Q:O QB:O VDDI:B VSSI:B
MM3 NET037 CKT VSSI VSSI nch_mac L=30N W=120N M=1
MM2 QB Q NET037 VSSI nch_mac L=30N W=120N M=1
MM11 QB IN NET38 VSSI nch_mac L=30N W=320N M=1
MM8 NET38 CKC VSSI VSSI nch_mac L=30N W=320N M=1
MM1 QB Q NET036 VDDI pch_mac L=30N W=120N M=1
MM0 NET036 CKC VDDI VDDI pch_mac L=30N W=120N M=1
MM9 NET39 CKT VDDI VDDI pch_mac L=30N W=430N M=1
MM10 QB IN NET39 VDDI pch_mac L=30N W=430N M=1
XI1 QB VSSI VSSI VDDI VDDI Q SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U MULTI=1 FP=1 
+ WP=0.43U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CNTWRAPER_LCH_M4_V3
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CNTWRAPER_LCH_M4_V3 AA[11] AA[10] AA[9] AA[8] AA[7] AA[6] AA[5] AA[4] 
+ AA[3] AA[2] AA[1] AA[0] AB[11] AB[10] AB[9] AB[8] AB[7] AB[6] AB[5] AB[4] 
+ AB[3] AB[2] AB[1] AB[0] AX[11] AX[10] AX[9] AX[8] AX[7] AX[6] AX[5] AX[4] 
+ AX[3] AX[2] AX[1] AX[0] CEBA CEBB CEBCA CEBCB CEBTA CEBTB CEX CEXBAF CKC CKT 
+ CLK DFF_SETB PHASESEL VDDI VSSI WEBA WEBB WEBCB WEBCBF WEBTB WEX
*.PININFO AA[11]:I AA[10]:I AA[9]:I AA[8]:I AA[7]:I AA[6]:I AA[5]:I AA[4]:I 
*.PININFO AA[3]:I AA[2]:I AA[1]:I AA[0]:I AB[11]:I AB[10]:I AB[9]:I AB[8]:I 
*.PININFO AB[7]:I AB[6]:I AB[5]:I AB[4]:I AB[3]:I AB[2]:I AB[1]:I AB[0]:I 
*.PININFO CEBA:I CEBB:I CKC:I CKT:I CLK:I DFF_SETB:I PHASESEL:I WEBA:I WEBB:I 
*.PININFO AX[11]:O AX[10]:O AX[9]:O AX[8]:O AX[7]:O AX[6]:O AX[5]:O AX[4]:O 
*.PININFO AX[3]:O AX[2]:O AX[1]:O AX[0]:O CEBCA:O CEBCB:O CEBTA:O CEBTB:O 
*.PININFO CEX:O CEXBAF:O WEBCB:O WEBCBF:O WEBTB:O WEX:O VDDI:B VSSI:B
XI32 PHASESEL VSSI VSSI VDDI VDDI SEL1B SDBM200W80_INV_BULK FN=5 WN=0.76U LN=0.03U 
+ MULTI=1 FP=5 WP=0.98U LP=0.03U
XCEB_LCHB CKC CKT CEBB CEBTB CEBCB VDDI VSSI SDBM200W80_LPLCH_CEB
XCEB_LCHA CKC CKT CEBA CEBTA CEBCA VDDI VSSI SDBM200W80_LPLCH_CEB
XA_MUX[11] AA[11] ABT[11] SEL1B PHASESEL AX[11] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[10] AA[10] ABT[10] SEL1B PHASESEL AX[10] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[9] AA[9] ABT[9] SEL1B PHASESEL AX[9] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[8] AA[8] ABT[8] SEL1B PHASESEL AX[8] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[7] AA[7] ABT[7] SEL1B PHASESEL AX[7] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[6] AA[6] ABT[6] SEL1B PHASESEL AX[6] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[5] AA[5] ABT[5] SEL1B PHASESEL AX[5] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[4] AA[4] ABT[4] SEL1B PHASESEL AX[4] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[3] AA[3] ABT[3] SEL1B PHASESEL AX[3] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[2] AA[2] ABT[2] SEL1B PHASESEL AX[2] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[1] AA[1] ABT[1] SEL1B PHASESEL AX[1] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_MUX[0] AA[0] ABT[0] SEL1B PHASESEL AX[0] VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XWEB_MUX WEBA WEBTB SEL1B PHASESEL WEX VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XCEB_MUX CEBA CEBTB SEL1B PHASESEL CEX VDDI VSSI SDBM200W80_PHASE_SEL_ADD_V1
XA_LCHB[11] CKC CKT AB[11] ABT[11] NET052[0] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[10] CKC CKT AB[10] ABT[10] NET052[1] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[9] CKC CKT AB[9] ABT[9] NET052[2] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[8] CKC CKT AB[8] ABT[8] NET052[3] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[7] CKC CKT AB[7] ABT[7] NET052[4] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[6] CKC CKT AB[6] ABT[6] NET052[5] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[5] CKC CKT AB[5] ABT[5] NET052[6] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[4] CKC CKT AB[4] ABT[4] NET052[7] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[3] CKC CKT AB[3] ABT[3] NET052[8] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[2] CKC CKT AB[2] ABT[2] NET052[9] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[1] CKC CKT AB[1] ABT[1] NET052[10] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XA_LCHB[0] CKC CKT AB[0] ABT[0] NET052[11] VDDI VSSI SDBM200W80_LPLCH_DE_ADD
XWEBB_LCH CKC CKT WEBB WEBTB WEBCB VDDI VSSI SDBM200W80_LPLCH_DE_ADD
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CNT_WP_M4_V5
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CNT_WP_M4_V5 AA[1] AA[0] AA[11] AA[10] AA[9] AA[8] AA[7] AA[6] AA[5] 
+ AA[4] AA[3] AA[2] AB[1] AB[0] AB[11] AB[10] AB[9] AB[8] AB[7] AB[6] AB[5] 
+ AB[4] AB[3] AB[2] AX[11] AX[10] AX[9] AX[8] AX[7] AX[6] AX[5] AX[4] AX[3] 
+ AX[2] AX[1] AX[0] CEBA CEBB CEX CKP1 CKP1_TRK CKP2 CKPB1 CKP_EN CKP_RSTB 
+ CKP_TRK CKT CLK CLKII CLKII_RED DCLK_L DCLK_R IOSAE PHASESEL_L PHASESEL_R 
+ PTSEL[0] PTSEL[1] QCLKBA_L QCLKBA_R QCLKBB_L QCLKBB_R REDEN TIE_H VDDI VSSI 
+ WEBA WEBB WEBX
*.PININFO AA[1]:I AA[0]:I AA[11]:I AA[10]:I AA[9]:I AA[8]:I AA[7]:I AA[6]:I 
*.PININFO AA[5]:I AA[4]:I AA[3]:I AA[2]:I AB[1]:I AB[0]:I AB[11]:I AB[10]:I 
*.PININFO AB[9]:I AB[8]:I AB[7]:I AB[6]:I AB[5]:I AB[4]:I AB[3]:I AB[2]:I 
*.PININFO CEBA:I CEBB:I CKP_RSTB:I CLK:I IOSAE:I PTSEL[0]:I PTSEL[1]:I REDEN:I 
*.PININFO TIE_H:I WEBA:I WEBB:I AX[11]:O AX[10]:O AX[9]:O AX[8]:O AX[7]:O 
*.PININFO AX[6]:O AX[5]:O AX[4]:O AX[3]:O AX[2]:O AX[1]:O AX[0]:O CEX:O CKP1:O 
*.PININFO CKP1_TRK:O CKP2:O CKPB1:O CKP_EN:O CKP_TRK:O CKT:O CLKII:O 
*.PININFO CLKII_RED:O DCLK_L:O DCLK_R:O PHASESEL_L:O PHASESEL_R:O QCLKBA_L:O 
*.PININFO QCLKBA_R:O QCLKBB_L:O QCLKBB_R:O WEBX:O VDDI:B VSSI:B
XI135 CKPB2 CKPB1 VSSI VSSI VDDI VDDI CLKII SDBM200W80_NAND_BULK FN1=3 WN1=1.2U 
+ LN1=0.03U FN2=3 WN2=1.2U LN2=0.03U FP2=2 WP2=1.2U LP2=0.03U MULTI=1 FP1=2 
+ WP1=1.2U LP1=0.03U
XI91 CKPB2 CKPB1 VSSI VSSI VDDI VDDI CLKII_RED SDBM200W80_NAND_BULK FN1=10 WN1=1.2U 
+ LN1=0.03U FN2=10 WN2=1.2U LN2=0.03U FP2=10 WP2=1.2U LP2=0.03U MULTI=1 FP1=10 
+ WP1=1.2U LP1=0.03U
XCLK_BUF CKC CKPB1_TRK CKPB_EN CKT VDDI VSSI DCLK_L DCLK_R SDBM200W80_CLK_BUF_DP_V2
XCKG CEAI CEBAI CEBBI CEBI CKP1 CKP2 PTSEL[0] PTSEL[1] CKPB1 CKPB1_TRK CKPB2 
+ CKPB_EN CKP_EN CKP_RSTB CKTA CLK TIE_H VDDI VSSI SDBM200W80_CKG_GEN_V7
MM45 CLKII_RED REDEN VSSI VSSI nch_mac L=30N W=1.2U M=4
MM44 VDDI REDEN VDDI VDDI pch_mac L=30N W=1.2U M=12
XCLK_QLATCH CEBAF CKPB1 CKPB2 CKP_RSTB CKTA CKTA2 IOSAE QCLKBA_L QCLKBA_R 
+ QCLKBB_L QCLKBB_R VDDI VSSI SDBM200W80_Q_LATCH_CLK_1007
XCNTPIN_WRCNT AA[11] AA[10] AA[9] AA[8] AA[7] AA[6] AA[5] AA[4] AA[3] AA[2] 
+ AA[1] AA[0] AB[11] AB[10] AB[9] AB[8] AB[7] AB[6] AB[5] AB[4] AB[3] AB[2] 
+ AB[1] AB[0] AX[11] AX[10] AX[9] AX[8] AX[7] AX[6] AX[5] AX[4] AX[3] AX[2] 
+ AX[1] AX[0] CEBA CEBB CEAI CEBI CEBAI CEBBI CEX CEBAF CKC CKT CLK CKPB2 
+ CKP_EN VDDI VSSI WEBA WEBB WEBI WEBCBF WEBBI WEBX SDBM200W80_CNTWRAPER_LCH_M4_V3
XI161 CKPB2 CKPB1_TRK CKPB1 VSSI VSSI VDDI VDDI CKP_TRK SDBM200W80_NAND3_BULK FN1=3 
+ WN1=0.76U LN1=0.03U FN2=3 WN2=0.76U LN2=0.03U FN3=3 WN3=0.76U LN3=0.03U 
+ FP3=1 WP3=0.32U LP3=0.03U FP2=3 WP2=0.43U LP2=0.03U MULTI=1 FP1=3 WP1=0.43U 
+ LP1=0.03U
XI154 NET022 VSSI VSSI VDDI VDDI NET071 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U 
+ MULTI=1 FP=1 WP=0.54U LP=0.03U
XI50 NET089 VSSI VSSI VDDI VDDI PHASESEL_L SDBM200W80_INV_BULK FN=4 WN=0.76U LN=0.03U 
+ MULTI=1 FP=4 WP=0.98U LP=0.03U
XI49 NET071 VSSI VSSI VDDI VDDI NET089 SDBM200W80_INV_BULK FN=1 WN=0.76U LN=0.03U 
+ MULTI=1 FP=1 WP=0.98U LP=0.03U
XI153 CKPB1_TRK VSSI VSSI VDDI VDDI CKP1_TRK SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U 
+ MULTI=1 FP=1 WP=0.43U LP=0.03U
XI152 CKP_EN VSSI VSSI VDDI VDDI NET022 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U 
+ MULTI=1 FP=1 WP=0.54U LP=0.03U
XI51 NET089 VSSI VSSI VDDI VDDI PHASESEL_R SDBM200W80_INV_BULK FN=4 WN=0.76U LN=0.03U 
+ MULTI=1 FP=4 WP=0.98U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    AWTD_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_AWTD_M4 AWT AWT2 VDDI VSSI
*.PININFO AWT:I AWT2:O VDDI:B VSSI:B
XINV1 AWT VSSI VSSI VDDI VDDI AWT1B SDBM200W80_INV_BULK FN=4 WN=430N LN=0.03U MULTI=1 
+ FP=6 WP=430N LP=0.03U
XINV0 AWT1B VSSI VSSI VDDI VDDI AWT2 SDBM200W80_INV_BULK FN=8 WN=0.76U LN=0.03U MULTI=1 
+ FP=12 WP=0.76U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    VHILO_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_VHILO_M4 VDDI VHI VLO VSSI
*.PININFO VHI:O VLO:O VDDI:B VSSI:B
MN3 VSSI Z2 Z1 VSSI nch_mac L=30N W=320N M=1
MN0 VSSI Z1 Z1 VSSI nch_mac L=30N W=320N M=1
MN1 VSSI Z2 VLO VSSI nch_mac L=30N W=0.76U M=4
MP7 Z2 Z1 VDDI VDDI pch_mac L=30N W=320N M=1
MP2 VHI Z1 VDDI VDDI pch_mac L=30N W=0.76U M=4
MP0 Z2 Z2 VDDI VDDI pch_mac L=30N W=320N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    TM_MODE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_TM_MODE CKP1 CKP2 TMA TMB TMB_EN TM_EN VDDI VSSI
*.PININFO CKP1:I CKP2:I TMA:I TMB:I TMB_EN:O TM_EN:O VDDI:B VSSI:B
XI638 TM_EN VSSI VSSI VDDI VDDI TMB_EN SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U 
+ MULTI=1 FP=1 WP=0.76U LP=0.03U
XI636 NET30 NET28 VSSI VSSI VDDI VDDI TM_EN SDBM200W80_NAND_BULK FN1=1 WN1=0.43U 
+ LN1=0.03U FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.76U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.76U LP1=0.03U
XI631 TMB CKP2 VSSI VSSI VDDI VDDI NET30 SDBM200W80_NAND_BULK FN1=1 WN1=0.43U LN1=0.03U 
+ FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.76U LP2=0.03U MULTI=1 FP1=1 WP1=0.76U 
+ LP1=0.03U
XI634 TMA CKP1 VSSI VSSI VDDI VDDI NET28 SDBM200W80_NAND_BULK FN1=1 WN1=0.43U LN1=0.03U 
+ FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.76U LP2=0.03U MULTI=1 FP1=1 WP1=0.76U 
+ LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    RESETD_TSEL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_RESETD_TSEL CKP V[0] V[1] VDDI VSSI TD_01_11 TD_10
*.PININFO CKP:I V[0]:I V[1]:I TD_01_11:O TD_10:O VDDI:B VSSI:B
MM0_MIXV_SSH Z4 NET37 VDDI VDDI pch_mac L=30N W=150N M=1
MM7_MIXV_SSH Z5 Z4 VDDI VDDI pch_mac L=30N W=150N M=1
MM31_MIXV_SSH NET37 CKP VDDI VDDI pch_mac L=30N W=150N M=1
MM3_MIXV_SSH Z4 NET37 VSSI VSSI nch_mac L=30N W=150N M=1
MM10_MIXV_SSH Z5 Z4 VSSI VSSI nch_mac L=30N W=150N M=1
MM22_MIXV_SSH NET37 CKP VSSI VSSI nch_mac L=30N W=150N M=1
XND5_MIXV_SSH Z5 V[1] VSSI VSSI VDDI VDDI TD_10 SDBM200W80_NAND_BULK FN1=1 WN1=0.32U 
+ LN1=0.03U FN2=1 WN2=0.32U LN2=0.03U FP2=1 WP2=0.23U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.23U LP1=0.03U
XND0_MIXV_SSH TD_10 CKP VSSI VSSI VDDI VDDI Z0 SDBM200W80_NAND_BULK FN1=1 WN1=0.43U 
+ LN1=0.03U FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.23U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.23U LP1=0.03U
XND1_MIXV_SSH V[0] Z0 VSSI VSSI VDDI VDDI TD_01_11 SDBM200W80_NAND_BULK FN1=1 WN1=0.87U 
+ LN1=0.03U FN2=1 WN2=0.87U LN2=0.03U FP2=1 WP2=0.65U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.65U LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    RESETD_TSEL_WT
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_RESETD_TSEL_WT CKPB VDDI VSSI OUT WV[0] WV[1]
*.PININFO CKPB:I WV[0]:I WV[1]:I OUT:O VDDI:B VSSI:B
XI90 Z5 WV[1] VSSI VSSI VDDI VDDI TD_10 SDBM200W80_NAND_BULK FN1=1 WN1=0.43U LN1=0.03U 
+ FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.32U LP2=0.03U MULTI=1 FP1=1 WP1=0.32U 
+ LP1=0.03U
XI97 TD_10 CKPB VSSI VSSI VDDI VDDI Z0 SDBM200W80_NAND_BULK FN1=1 WN1=0.43U LN1=0.03U 
+ FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.32U LP2=0.03U MULTI=1 FP1=1 WP1=0.32U 
+ LP1=0.03U
XI98 WV[0] Z0 VSSI VSSI VDDI VDDI TD_01_11 SDBM200W80_NAND_BULK FN1=1 WN1=0.43U 
+ LN1=0.03U FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.32U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.32U LP1=0.03U
XI87_MIXV_SLH TD_10 TD_01_11 VSSI VSSI VDDI VDDI NET78 SDBM200W80_NAND_BULK FN1=1 
+ WN1=0.43U LN1=0.03U FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.32U LP2=0.03U 
+ MULTI=1 FP1=1 WP1=0.32U LP1=0.03U
XI95 Z4 VSSI VSSI VDDI VDDI Z5 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 FP=1 
+ WP=0.15U LP=0.03U
XI93 Z3 VSSI VSSI VDDI VDDI Z4 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 FP=1 
+ WP=0.15U LP=0.03U
XI91 CKPB VSSI VSSI VDDI VDDI Z3 SDBM200W80_INV_BULK FN=1 WN=0.15U LN=0.03U MULTI=1 
+ FP=1 WP=0.15U LP=0.03U
XI89_MIXV_SLH NET78 VSSI VSSI VDDI VDDI OUT SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.32U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DECB1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DECB1 CKP CLK DEC PREDEC VDDI VSSI
*.PININFO CKP:I CLK:I PREDEC:I DEC:O VDDI:B VSSI:B
MTN1 NT1 CKP NT3 VSSI nch_mac L=30N W=430N M=1
MTN2 NT3 PREDEC VSSI VSSI nch_mac L=30N W=0.74U M=5
MM0 NT1 CLK NT3 VSSI nch_mac L=30N W=0.74U M=3
MN0 DEC NT1 VSSI VSSI nch_mac L=30N W=0.74U M=6
MM8 NT1 CKP NET31 VDDI pch_mac L=30N W=0.64U M=2
MM1 NET31 CLK VDDI VDDI pch_mac L=30N W=0.64U M=2
MM3 NT1 PREDEC VDDI VDDI pch_mac L=30N W=430N M=1
MP0 DEC NT1 VDDI VDDI pch_mac L=30N W=0.74U M=12
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DEC_Y
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DEC_Y CKP CLK DEC PREDEC VDDI VSSI
*.PININFO CKP:I CLK:I PREDEC:I DEC:O VDDI:B VSSI:B
MTN1 NT1 CKP NT3 VSSI nch_mac L=30N W=430N M=1
MTN2 NT3 PREDEC VSSI VSSI nch_mac L=30N W=0.74U M=5
MM0 NT1 CLK NT3 VSSI nch_mac L=30N W=0.74U M=3
MN0 DEC NT1 VSSI VSSI nch_mac L=30N W=0.74U M=6
MM1 NET31 CLK VDDI VDDI pch_mac L=30N W=0.64U M=2
MM8 NT1 CKP NET31 VDDI pch_mac L=30N W=0.64U M=2
MM3 NT1 PREDEC VDDI VDDI pch_mac L=30N W=430N M=1
MP0 DEC NT1 VDDI VDDI pch_mac L=30N W=0.74U M=12
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DECB4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DECB4 IN0A IN0B IN1A IN1B IN2 PREDEC0 PREDEC1 PREDEC2 PREDEC3 VDDI VSSI
*.PININFO IN0A:I IN0B:I IN1A:I IN1B:I IN2:I PREDEC0:O PREDEC1:O PREDEC2:O 
*.PININFO PREDEC3:O VDDI:B VSSI:B
MM19 N5 IN1B NET19 VSSI nch_mac L=30N W=430N M=1
MM20 NET0154 IN0B N5 VSSI nch_mac L=30N W=300N M=1
MM21 NET0150 IN0A N5 VSSI nch_mac L=30N W=300N M=1
MM26 NET19 IN2 VSSI VSSI nch_mac L=30N W=430N M=2
MM8 N2 IN1A NET19 VSSI nch_mac L=30N W=430N M=1
MM7 NET0138 IN0B N2 VSSI nch_mac L=30N W=300N M=1
MM0 NET0134 IN0A N2 VSSI nch_mac L=30N W=300N M=1
MM15 NET0154 IN1B VDDI VDDI pch_mac L=30N W=250N M=1
MM16 NET0154 IN0B VDDI VDDI pch_mac L=30N W=250N M=1
MM17 NET0150 IN1B VDDI VDDI pch_mac L=30N W=250N M=1
MM18 NET0150 IN0A VDDI VDDI pch_mac L=30N W=250N M=1
MM22 NET0150 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM23 NET0154 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM24 NET0138 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM25 NET0134 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM5 NET0138 IN1A VDDI VDDI pch_mac L=30N W=250N M=1
MM4 NET0138 IN0B VDDI VDDI pch_mac L=30N W=250N M=1
MM2 NET0134 IN1A VDDI VDDI pch_mac L=30N W=250N M=1
MM1 NET0134 IN0A VDDI VDDI pch_mac L=30N W=250N M=1
XINV3 NET0154 VSSI VSSI VDDI VDDI PREDEC3 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV2 NET0150 VSSI VSSI VDDI VDDI PREDEC2 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV1 NET0138 VSSI VSSI VDDI VDDI PREDEC1 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV0 NET0134 VSSI VSSI VDDI VDDI PREDEC0 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DECB1_DCLK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DECB1_DCLK CKPDCLK CLK DEC PREDEC VDDI VSSI
*.PININFO CKPDCLK:I CLK:I PREDEC:I DEC:O VDDI:B VSSI:B
MM0 NT1 CLK NT3 VSSI nch_mac L=30N W=0.74U M=3
MN0 DEC NT1 VSSI VSSI nch_mac L=30N W=0.74U M=10
MTN1 NT1 CKPDCLK NT3 VSSI nch_mac L=30N W=430N M=1
MTN2 NT3 PREDEC VSSI VSSI nch_mac L=30N W=0.74U M=5
MM2 NT1 CKPDCLK NET59 VDDI pch_mac L=30N W=0.74U M=2
MM1 NET59 CLK VDDI VDDI pch_mac L=30N W=0.74U M=2
MM3 NT1 PREDEC VDDI VDDI pch_mac L=30N W=430N M=1
MP0 DEC NT1 VDDI VDDI pch_mac L=30N W=0.74U M=12
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    ABUF_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_ABUF_WOBIST A AC AT AX1B CK1B CK2 VDDI VSSI
*.PININFO A:I CK1B:I CK2:I AC:O AT:O AX1B:O VDDI:B VSSI:B
MM23 NET0108 CK1B VSSI VSSI nch_mac L=30N W=380N M=2
MM21 NET078 AC VSSI VSSI nch_mac L=30N W=120N M=1
MM20 AT CK2 NET078 VSSI nch_mac L=30N W=120N M=1
MM19 AT A NET0108 VSSI nch_mac L=30N W=380N M=2
MM29 AT A NET0145 VDDI pch_mac L=30N W=0.54U M=2
MM28 NET0145 CK2 VDDI VDDI pch_mac L=30N W=0.54U M=2
MM27 NET0149 AC VDDI VDDI pch_mac L=30N W=120N M=1
MM26 AT CK1B NET0149 VDDI pch_mac L=30N W=120N M=1
XI25 AT VSSI VSSI VDDI VDDI AC SDBM200W80_INV_BULK FN=2 WN=0.4U LN=0.03U MULTI=1 FP=2 
+ WP=0.52U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    ABUF_DECB4_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_ABUF_DECB4_WOBIST CK1B CK2 IN[0] IN[1] IN[2] OUT[0] OUT[1] OUT[2] 
+ OUT[3] OUT[4] OUT[5] OUT[6] OUT[7] VDDI VSSI
*.PININFO CK1B:I CK2:I IN[0]:I IN[1]:I IN[2]:I OUT[0]:O OUT[1]:O OUT[2]:O 
*.PININFO OUT[3]:O OUT[4]:O OUT[5]:O OUT[6]:O OUT[7]:O VDDI:B VSSI:B
XABUF[2] IN[2] AXC[2] AXT[2] AX[2] CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XABUF[1] IN[1] AXC[1] AXT[1] AX[1] CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XABUF[0] IN[0] AXC[0] AXT[0] AX[0] CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XDECB4[0] AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] OUT[0] OUT[1] OUT[2] OUT[3] VDDI 
+ VSSI SDBM200W80_DECB4
XDECB4[1] AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] OUT[4] OUT[5] OUT[6] OUT[7] VDDI 
+ VSSI SDBM200W80_DECB4
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    ABUF_WEB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_ABUF_WEB A AC AT AX1B CK1B CK2 VDDI VSSI
*.PININFO A:I CK1B:I CK2:I AC:O AT:O AX1B:O VDDI:B VSSI:B
MM23 NET0108 CK1B VSSI VSSI nch_mac L=30N W=380N M=2
MM21 NET078 AC VSSI VSSI nch_mac L=30N W=120N M=1
MM20 AT CK2 NET078 VSSI nch_mac L=30N W=120N M=1
MM19 AT A NET0108 VSSI nch_mac L=30N W=380N M=2
MM29 AT A NET0145 VDDI pch_mac L=30N W=320N M=2
MM28 NET0145 CK2 VDDI VDDI pch_mac L=30N W=320N M=2
MM27 NET0149 AC VDDI VDDI pch_mac L=30N W=120N M=1
MM26 AT CK1B NET0149 VDDI pch_mac L=30N W=120N M=1
XI25 AT VSSI VSSI VDDI VDDI AC SDBM200W80_INV_BULK FN=2 WN=0.4U LN=0.03U MULTI=1 FP=2 
+ WP=0.52U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DECB1_DCLKA
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DECB1_DCLKA CKPDCLK CLK DEC PREDEC VDDI VSSI
*.PININFO CKPDCLK:I CLK:I PREDEC:I DEC:O VDDI:B VSSI:B
MM0 NT1 CLK NT3 VSSI nch_mac L=30N W=0.74U M=3
MN0 DEC NT1 VSSI VSSI nch_mac L=30N W=0.8U M=6
MTN1 NT1 CKPDCLK NT3 VSSI nch_mac L=30N W=430N M=1
MTN2 NT3 PREDEC VSSI VSSI nch_mac L=30N W=0.74U M=5
MM2 NT1 CKPDCLK NET59 VDDI pch_mac L=30N W=0.65U M=2
MM1 NET59 CLK VDDI VDDI pch_mac L=30N W=0.65U M=2
MM3 NT1 PREDEC VDDI VDDI pch_mac L=30N W=430N M=1
MP0 DEC NT1 VDDI VDDI pch_mac L=30N W=0.74U M=12
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DECB1_BS_SEG
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DECB1_BS_SEG CKP CLK DEC PREDEC VDDI VSSI
*.PININFO CKP:I CLK:I PREDEC:I DEC:O VDDI:B VSSI:B
MM3 NT1 PREDEC VDDI VDDI pch_mac L=30N W=430N M=1
MP0 DEC NT1 VDDI VDDI pch_mac L=30N W=0.74U M=12
MM1 NT1 CLK VDDI VDDI pch_mac L=30N W=0.64U M=2
MTN1 NT1 CLK NT3 VSSI nch_mac L=30N W=430N M=1
MTN2 NT3 PREDEC VSSI VSSI nch_mac L=30N W=0.74U M=5
MM0 NT1 CLK NT3 VSSI nch_mac L=30N W=0.74U M=3
MN0 DEC NT1 VSSI VSSI nch_mac L=30N W=0.74U M=7
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DECB4_Y
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DECB4_Y IN0A IN0B IN1A IN1B IN2 PREDEC0 PREDEC1 PREDEC2 PREDEC3 VDDI 
+ VSSI
*.PININFO IN0A:I IN0B:I IN1A:I IN1B:I IN2:I PREDEC0:O PREDEC1:O PREDEC2:O 
*.PININFO PREDEC3:O VDDI:B VSSI:B
MM19 N5 IN1B NET19 VSSI nch_mac L=30N W=430N M=1
MM20 NET0154 IN0B N5 VSSI nch_mac L=30N W=300N M=1
MM21 NET0150 IN0A N5 VSSI nch_mac L=30N W=300N M=1
MM26 NET19 IN2 VSSI VSSI nch_mac L=30N W=280N M=2
MM8 N2 IN1A NET19 VSSI nch_mac L=30N W=430N M=1
MM7 NET0138 IN0B N2 VSSI nch_mac L=30N W=300N M=1
MM0 NET0134 IN0A N2 VSSI nch_mac L=30N W=300N M=1
MM15 NET0154 IN1B VDDI VDDI pch_mac L=30N W=250N M=1
MM16 NET0154 IN0B VDDI VDDI pch_mac L=30N W=250N M=1
MM17 NET0150 IN1B VDDI VDDI pch_mac L=30N W=250N M=1
MM18 NET0150 IN0A VDDI VDDI pch_mac L=30N W=250N M=1
MM22 NET0150 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM23 NET0154 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM24 NET0138 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM25 NET0134 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM5 NET0138 IN1A VDDI VDDI pch_mac L=30N W=250N M=1
MM4 NET0138 IN0B VDDI VDDI pch_mac L=30N W=250N M=1
MM2 NET0134 IN1A VDDI VDDI pch_mac L=30N W=250N M=1
MM1 NET0134 IN0A VDDI VDDI pch_mac L=30N W=250N M=1
XINV3 NET0154 VSSI VSSI VDDI VDDI PREDEC3 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV2 NET0150 VSSI VSSI VDDI VDDI PREDEC2 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV1 NET0138 VSSI VSSI VDDI VDDI PREDEC1 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV0 NET0134 VSSI VSSI VDDI VDDI PREDEC0 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    DECB4_Z0
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_DECB4_Z0 IN0A IN0B IN1A IN1B IN2 PREDEC0 PREDEC1 PREDEC2 PREDEC3 VDDI 
+ VSSI
*.PININFO IN0A:I IN0B:I IN1A:I IN1B:I IN2:I PREDEC0:O PREDEC1:O PREDEC2:O 
*.PININFO PREDEC3:O VDDI:B VSSI:B
MM19 N5 IN1B NET19 VSSI nch_mac L=30N W=430N M=1
MM20 NET0154 IN0B N5 VSSI nch_mac L=30N W=300N M=1
MM21 NET0150 IN0A N5 VSSI nch_mac L=30N W=300N M=1
MM26 NET19 IN2 VSSI VSSI nch_mac L=30N W=430N M=2
MM8 N2 IN1A NET19 VSSI nch_mac L=30N W=430N M=1
MM7 NET0138 IN0B N2 VSSI nch_mac L=30N W=300N M=1
MM0 NET0134 IN0A N2 VSSI nch_mac L=30N W=300N M=1
MM15 NET0154 IN1B VDDI VDDI pch_mac L=30N W=250N M=1
MM16 NET0154 IN0B VDDI VDDI pch_mac L=30N W=250N M=1
MM17 NET0150 IN1B VDDI VDDI pch_mac L=30N W=250N M=1
MM18 NET0150 IN0A VDDI VDDI pch_mac L=30N W=250N M=1
MM22 NET0150 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM23 NET0154 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM24 NET0138 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM25 NET0134 IN2 VDDI VDDI pch_mac L=30N W=250N M=1
MM5 NET0138 IN1A VDDI VDDI pch_mac L=30N W=250N M=1
MM4 NET0138 IN0B VDDI VDDI pch_mac L=30N W=250N M=1
MM2 NET0134 IN1A VDDI VDDI pch_mac L=30N W=250N M=1
MM1 NET0134 IN0A VDDI VDDI pch_mac L=30N W=250N M=1
XINV3 NET0154 VSSI VSSI VDDI VDDI PREDEC3 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV2 NET0150 VSSI VSSI VDDI VDDI PREDEC2 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV1 NET0138 VSSI VSSI VDDI VDDI PREDEC1 SDBM200W80_INV_BULK FN=1 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
XINV0 NET0134 VSSI VSSI VDDI VDDI PREDEC0 SDBM200W80_INV_BULK FN=2 WN=0.30U LN=0.03U 
+ MULTI=1 FP=2 WP=0.30U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    ABUF_DECB4_WOBIST_Z0
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_ABUF_DECB4_WOBIST_Z0 CK1B CK2 IN[0] IN[1] IN[2] OUT[0] OUT[1] OUT[2] 
+ OUT[3] OUT[4] OUT[5] OUT[6] OUT[7] VDDI VSSI
*.PININFO CK1B:I CK2:I IN[0]:I IN[1]:I IN[2]:I OUT[0]:O OUT[1]:O OUT[2]:O 
*.PININFO OUT[3]:O OUT[4]:O OUT[5]:O OUT[6]:O OUT[7]:O VDDI:B VSSI:B
XABUF[2] IN[2] AXC[2] AXT[2] AX[2] CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XABUF[1] IN[1] AXC[1] AXT[1] AX[1] CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XABUF[0] IN[0] AXC[0] AXT[0] AX[0] CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XDECB4[1] AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] OUT[4] OUT[5] OUT[6] OUT[7] VDDI 
+ VSSI SDBM200W80_DECB4
XDECB4[0] AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] OUT[0] OUT[1] OUT[2] OUT[3] VDDI 
+ VSSI SDBM200W80_DECB4_Z0
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CDEC_M4_WOBIST_RED_DP_V4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CDEC_M4_WOBIST_RED_DP_V4 CEB CK1B CK2 CK2_TRK CKD CKP CKPD CKPDCLK 
+ CKPD_RED CKP_RED DCLKA DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ REDEN VDDI VSSI WEB WEB2 WEB5B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] Y[0] Y[1]
*.PININFO CEB:I CK1B:I CK2:I CK2_TRK:I CKP:I CKPD:I CKPDCLK:I CKPD_RED:I 
*.PININFO CKP_RED:I REDEN:I WEB:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I 
*.PININFO X[6]:I X[7]:I X[8]:I X[9]:I Y[0]:I Y[1]:I CKD:O DCLKA:O DEC_X0[0]:O 
*.PININFO DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O 
*.PININFO DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O 
*.PININFO DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O 
*.PININFO DEC_X2[0]:O DEC_X2[1]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O 
*.PININFO DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O 
*.PININFO DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O 
*.PININFO DEC_Y[6]:O DEC_Y[7]:O WEB2:O WEB5B:O VDDI:B VSSI:B
XIDEC_X2[0] CKPD_RED CKP_RED DEC_X2[0] XC[0] VDDI VSSI SDBM200W80_DECB1
XIDEC_X2[1] CKPD_RED CKP_RED DEC_X2[1] XC[1] VDDI VSSI SDBM200W80_DECB1
XIDEC_X0[0] CKPD_RED CKP_RED DEC_X0[0] XA[0] VDDI VSSI SDBM200W80_DECB1
XIDEC_X0[1] CKPD_RED CKP_RED DEC_X0[1] XA[1] VDDI VSSI SDBM200W80_DECB1
XIDEC_X0[2] CKPD_RED CKP_RED DEC_X0[2] XA[2] VDDI VSSI SDBM200W80_DECB1
XIDEC_X0[3] CKPD_RED CKP_RED DEC_X0[3] XA[3] VDDI VSSI SDBM200W80_DECB1
XIDEC_X0[4] CKPD_RED CKP_RED DEC_X0[4] XA[4] VDDI VSSI SDBM200W80_DECB1
XIDEC_X0[5] CKPD_RED CKP_RED DEC_X0[5] XA[5] VDDI VSSI SDBM200W80_DECB1
XIDEC_X0[6] CKPD_RED CKP_RED DEC_X0[6] XA[6] VDDI VSSI SDBM200W80_DECB1
XIDEC_X0[7] CKPD_RED CKP_RED DEC_X0[7] XA[7] VDDI VSSI SDBM200W80_DECB1
XIDEC_X1[0] CKPD_RED CKP_RED DEC_X1[0] XB[0] VDDI VSSI SDBM200W80_DECB1
XIDEC_X1[1] CKPD_RED CKP_RED DEC_X1[1] XB[1] VDDI VSSI SDBM200W80_DECB1
XIDEC_X1[2] CKPD_RED CKP_RED DEC_X1[2] XB[2] VDDI VSSI SDBM200W80_DECB1
XIDEC_X1[3] CKPD_RED CKP_RED DEC_X1[3] XB[3] VDDI VSSI SDBM200W80_DECB1
XIDEC_X1[4] CKPD_RED CKP_RED DEC_X1[4] XB[4] VDDI VSSI SDBM200W80_DECB1
XIDEC_X1[5] CKPD_RED CKP_RED DEC_X1[5] XB[5] VDDI VSSI SDBM200W80_DECB1
XIDEC_X1[6] CKPD_RED CKP_RED DEC_X1[6] XB[6] VDDI VSSI SDBM200W80_DECB1
XIDEC_X1[7] CKPD_RED CKP_RED DEC_X1[7] XB[7] VDDI VSSI SDBM200W80_DECB1
XIDEC_Y[0] CKPD CKP DEC_Y[0] XY[0] VDDI VSSI SDBM200W80_DEC_Y
XIDEC_Y[1] CKPD CKP DEC_Y[1] XY[1] VDDI VSSI SDBM200W80_DEC_Y
XIDEC_Y[2] CKPD CKP DEC_Y[2] XY[2] VDDI VSSI SDBM200W80_DEC_Y
XIDEC_Y[3] CKPD CKP DEC_Y[3] XY[3] VDDI VSSI SDBM200W80_DEC_Y
XIDEC_Y[4] CKPD CKP DEC_Y[4] XY[4] VDDI VSSI SDBM200W80_DEC_Y
XIDEC_Y[5] CKPD CKP DEC_Y[5] XY[5] VDDI VSSI SDBM200W80_DEC_Y
XIDEC_Y[6] CKPD CKP DEC_Y[6] XY[6] VDDI VSSI SDBM200W80_DEC_Y
XIDEC_Y[7] CKPD CKP DEC_Y[7] XY[7] VDDI VSSI SDBM200W80_DEC_Y
XI345 NET051 VSSI VSSI VDDI VDDI XC[1] SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U 
+ MULTI=1 FP=1 WP=0.6U LP=0.03U
XI347 WEB3B VSSI VSSI VDDI VDDI NET044 SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U 
+ MULTI=1 FP=1 WP=0.43U LP=0.03U
XI348 NET044 VSSI VSSI VDDI VDDI NET023 SDBM200W80_INV_BULK FN=2 WN=0.43U LN=0.03U 
+ MULTI=1 FP=2 WP=0.65U LP=0.03U
XI354 CK1B VSSI VSSI VDDI VDDI CKP1D SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.43U LP=0.03U
XI355 CK2_TRK VSSI VSSI VDDI VDDI CK1B_TRK SDBM200W80_INV_BULK FN=1 WN=0.32U LN=0.03U 
+ MULTI=1 FP=1 WP=0.43U LP=0.03U
XI356 WEB VSSI VSSI VDDI VDDI NET019 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U MULTI=1 
+ FP=1 WP=0.32U LP=0.03U
XINV0 REDEN VSSI VSSI VDDI VDDI NET30 SDBM200W80_INV_BULK FN=1 WN=0.27U LN=0.03U 
+ MULTI=1 FP=1 WP=0.54U LP=0.03U
XI350 XC[1] VSSI VSSI VDDI VDDI XC[0] SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U 
+ MULTI=1 FP=1 WP=0.6U LP=0.03U
XIPDEC_Y[1] AYC[0] AYT[0] AYC[1] AYT[1] WEB3B XY[4] XY[5] XY[6] XY[7] VDDI 
+ VSSI SDBM200W80_DECB4
XIDEC_CKD CKPD CKP CKD NET023 VDDI VSSI SDBM200W80_DECB1_DCLK
MM13 Z[0] NET30 Z0_REDEN VSSI nch_mac L=30N W=540N M=1
XABUF_PDEC_X0 CK1B CK2 X[0] X[1] X[2] XA[0] XA[1] XA[2] XA[3] XA[4] XA[5] 
+ XA[6] XA[7] VDDI VSSI SDBM200W80_ABUF_DECB4_WOBIST
XABUF_PDEC_X1 CK1B CK2 X[3] X[4] X[5] XB[0] XB[1] XB[2] XB[3] XB[4] XB[5] 
+ XB[6] XB[7] VDDI VSSI SDBM200W80_ABUF_DECB4_WOBIST
XWEBBUF WEB WEB3B WEB2 NET032 CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WEB
MM0 Z0_REDEN NET30 VDDI VDDI pch_mac L=30N W=540N M=1
MM12 Z[0] REDEN Z0_REDEN VDDI pch_mac L=30N W=540N M=1
XIDEC_DCLKA CKP1D CK2 DCLKA NET023 VDDI VSSI SDBM200W80_DECB1_DCLKA
XIDEC_X3[1] CKPD_RED CKP_RED DEC_X3[1] Z[1] VDDI VSSI SDBM200W80_DECB1_BS_SEG
XIDEC_X3[2] CKPD_RED CKP_RED DEC_X3[2] Z[2] VDDI VSSI SDBM200W80_DECB1_BS_SEG
XIDEC_X3[3] CKPD_RED CKP_RED DEC_X3[3] Z[3] VDDI VSSI SDBM200W80_DECB1_BS_SEG
XIDEC_X3[4] CKPD_RED CKP_RED DEC_X3[4] Z[4] VDDI VSSI SDBM200W80_DECB1_BS_SEG
XIDEC_X3[5] CKPD_RED CKP_RED DEC_X3[5] Z[5] VDDI VSSI SDBM200W80_DECB1_BS_SEG
XIDEC_X3[6] CKPD_RED CKP_RED DEC_X3[6] Z[6] VDDI VSSI SDBM200W80_DECB1_BS_SEG
XIDEC_X3[7] CKPD_RED CKP_RED DEC_X3[7] Z[7] VDDI VSSI SDBM200W80_DECB1_BS_SEG
XIDEC_X3[0] CKP CKP DEC_X3[0] Z0_REDEN VDDI VSSI SDBM200W80_DECB1_BS_SEG
XI338 CEB NET019 VSSI VSSI VDDI VDDI NET045 SDBM200W80_NAND_BULK FN1=1 WN1=0.43U 
+ LN1=0.03U FN2=1 WN2=0.43U LN2=0.03U FP2=1 WP2=0.21U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.21U LP1=0.03U
XI352 NET045 WEB5B CEB2 NET038 CK1B_TRK CK2_TRK VDDI VSSI SDBM200W80_ABUF_WOBIST
XI343[0] X[6] NET051 NET034 NET036 CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XABUF_Y[0] Y[0] AYC[0] AYT[0] AY[0] CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XABUF_Y[1] Y[1] AYC[1] AYT[1] AY[1] CK1B CK2 VDDI VSSI SDBM200W80_ABUF_WOBIST
XIPDEC_Y[0] AYC[0] AYT[0] AYC[1] AYT[1] WEB2 XY[0] XY[1] XY[2] XY[3] VDDI VSSI 
+ SDBM200W80_DECB4_Y
XABUF_PDEC_X3 CK1B CK2 X[7] X[8] X[9] Z[0] Z[1] Z[2] Z[3] Z[4] Z[5] Z[6] Z[7] 
+ VDDI VSSI SDBM200W80_ABUF_DECB4_WOBIST_Z0
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    RESETD_M4_RED_DP_V3_H
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_RESETD_M4_RED_DP_V3_H BLTRKWLDRV CKP CKP1 CKP2 CKPD CKPDCLK CKPD_RED 
+ CKP_RED CKP_TRK CLK IOSAEB QLATCH RSC RSC_TRK_H RSC_TRK_W TMA TMB TRKBL VDDI 
+ VSSI WEBXL WLP_SAE WLP_SAE_TK RV[0] RV[1] WV[0] WV[1]
*.PININFO CKP:I CKP1:I CKP2:I CKP_RED:I CKP_TRK:I CLK:I TMA:I TMB:I WEBXL:I 
*.PININFO RV[0]:I RV[1]:I WV[0]:I WV[1]:I BLTRKWLDRV:O CKPD:O CKPDCLK:O 
*.PININFO CKPD_RED:O IOSAEB:O QLATCH:O RSC:O WLP_SAE:O RSC_TRK_H:B RSC_TRK_W:B 
*.PININFO TRKBL:B VDDI:B VSSI:B WLP_SAE_TK:B
XI649 CKP1 CKP2 TMA TMB TMB_EN TM_EN VDDI VSSI SDBM200W80_TM_MODE
MM28 NET0310 TRKBL1B VDDI VDDI pch_mac L=30N W=320N M=1
MM33_MIXV_SSH NET0256 NET0215 NET0293 VDDI pch_mac L=30N W=150N M=1
MM32_MIXV_SSH NET0215 NET0206 VDDI VDDI pch_mac L=30N W=150N M=1
MM10 TRKBL1B TRKBL NET0298 VDDI pch_mac L=30N W=980N M=1
MM12 NET0298 TM_EN VDDI VDDI pch_mac L=30N W=0.98U M=3
MM16_MIXV_SSH NET0206 WLP_SAE NET0295 VDDI pch_mac L=30N W=150N M=1
MM34_MIXV_SSH NET0293 NET0215 VDDI VDDI pch_mac L=30N W=150N M=1
MM15_MIXV_SSH NET0295 WLP_SAE VDDI VDDI pch_mac L=30N W=150N M=1
MM27 NET0311 D7 VDDI VDDI pch_mac L=30N W=120N M=1
MM29 AXL WEBXL NET0310 VDDI pch_mac L=30N W=320N M=1
MM26 AXL TRKBL2B NET0311 VDDI pch_mac L=30N W=120N M=1
MP16 WLP_SAE TRKBL2 VDDI VDDI pch_mac L=30N W=1.2U M=13
MM30 NET0299 TMB_EN VDDI VDDI pch_mac L=30N W=430N M=1
MM8 TRKBL1B NET0147 NET0299 VDDI pch_mac L=30N W=430N M=1
XI637 TRKBL_TM CLK_TM VSSI VSSI VDDI VDDI NET0147 SDBM200W80_NAND_BULK FN1=1 WN1=0.43U 
+ LN1=30N FN2=1 WN2=0.43U LN2=30N FP2=1 WP2=0.21U LP2=30N MULTI=1 FP1=1 
+ WP1=0.21U LP1=30N
XI521 TRKBL2 WLP_SAE_TK1B VSSI VSSI VDDI VDDI QLATCH SDBM200W80_NAND_BULK FN1=2 
+ WN1=1.2U LN1=0.03U FN2=2 WN2=1.2U LN2=0.03U FP2=1 WP2=0.76U LP2=0.03U 
+ MULTI=1 FP1=3 WP1=1.15U LP1=0.03U
XI574_MIXV_SLH NET0194 TRKBL1B VSSI VSSI VDDI VDDI RSTCKB SDBM200W80_NAND_BULK FN1=1 
+ WN1=0.98U LN1=30N FN2=1 WN2=0.98U LN2=30N FP2=1 WP2=540N LP2=30N MULTI=1 
+ FP1=1 WP1=540N LP1=30N
XI624 CKP_TRK RV[0] RV[1] VDDI VSSI RTD_01_11 RTD_10 SDBM200W80_RESETD_TSEL
XI665 RSC_TRK_H RSC_TRK_W VSSI VSSI VDDI VDDI Z8_TRK SDBM200W80_NOR_BULK FN1=2 
+ WN1=0.56U LN1=0.03U FN2=2 WN2=0.56U LN2=0.03U FP2=2 WP2=0.56U LP2=0.03U 
+ MULTI=1 FP1=2 WP1=0.56U LP1=0.03U
XNOR0 Z8_TRK RSTCKB VSSI VSSI VDDI VDDI RSTCK SDBM200W80_NOR_BULK FN1=2 WN1=0.76U 
+ LN1=0.03U FN2=2 WN2=0.76U LN2=0.03U FP2=2 WP2=1.2U LP2=0.03U MULTI=1 FP1=2 
+ WP1=1.2U LP1=0.03U
XI625_MIXV_SLH D7 TRKBL2B VSSI VSSI VDDI VDDI TRKBL3B SDBM200W80_NOR_BULK FN1=1 
+ WN1=0.76U LN1=0.03U FN2=2 WN2=0.76U LN2=0.03U FP2=2 WP2=0.98U LP2=0.03U 
+ MULTI=1 FP1=3 WP1=0.98U LP1=0.03U
MM9 NET0297 TMB_EN VSSI VSSI nch_mac L=30N W=0.65U M=3
MM43_MIXV_SSH NET0215 NET0206 NET0294 VSSI nch_mac L=30N W=150N M=1
MM21 NET0308 D7 VSSI VSSI nch_mac L=30N W=120N M=1
MM19 AXL WEBXL NET0296 VSSI nch_mac L=30N W=210N M=1
MM46_MIXV_SSH NET0256 NET0215 VSSI VSSI nch_mac L=30N W=150N M=1
MM1 TRKBL1B NET0147 NET0300 VSSI nch_mac L=30N W=540N M=1
MM2 NET0300 TM_EN VSSI VSSI nch_mac L=30N W=540N M=1
MM44_MIXV_SSH NET0294 NET0206 VSSI VSSI nch_mac L=30N W=150N M=1
MN7 WLP_SAE TRKBL2 VSSI VSSI nch_mac L=30N W=1.2U M=7
MM18_MIXV_SSH NET0206 WLP_SAE VSSI VSSI nch_mac L=30N W=150N M=1
MM20 AXL TRKBL1B NET0308 VSSI nch_mac L=30N W=120N M=1
MM23 NET0296 TRKBL2B VSSI VSSI nch_mac L=30N W=210N M=1
MM11 TRKBL1B TRKBL NET0297 VSSI nch_mac L=30N W=650N M=1
XI664 NET0108 VSSI VSSI VDDI VDDI RSC_TRK_H SDBM200W80_INV_BULK FN=4 WN=0.8U LN=0.03U 
+ MULTI=1 FP=4 WP=1.2U LP=0.03U
XI618_MIXV_SLH TRKBL1B VSSI VSSI VDDI VDDI TRKBL2B SDBM200W80_INV_BULK FN=1 WN=0.98U 
+ LN=30N MULTI=1 FP=1 WP=1.09U LP=30N
XI633 RSTCK VSSI VSSI VDDI VDDI RSC SDBM200W80_INV_BULK FN=4 WN=0.87U LN=30N MULTI=1 
+ FP=4 WP=1.2U LP=30N
XI626_MIXV_SLH TRKBL3B VSSI VSSI VDDI VDDI TRKBL2 SDBM200W80_INV_BULK FN=3 WN=0.98U 
+ LN=30N MULTI=1 FP=3 WP=1.2U LP=30N
XI566 WLP_SAE_TK VSSI VSSI VDDI VDDI WLP_SAE_TK1B SDBM200W80_INV_BULK FN=1 WN=1.2U 
+ LN=0.03U MULTI=1 FP=1 WP=1.2U LP=0.03U
XI532 NET096 VSSI VSSI VDDI VDDI IOSAEB SDBM200W80_INV_BULK FN=8 WN=0.87U LN=0.03U 
+ MULTI=1 FP=8 WP=1.2U LP=0.03U
XI537 RTKB VSSI VSSI VDDI VDDI BLTRKWLDRV SDBM200W80_INV_BULK FN=9 WN=650N LN=30N 
+ MULTI=1 FP=9 WP=980N LP=30N
XI639 CLK VSSI VSSI VDDI VDDI CLK_TM SDBM200W80_INV_BULK FN=1 WN=0.12U LN=30N MULTI=1 
+ FP=1 WP=0.21U LP=30N
XI663 NET0108 VSSI VSSI VDDI VDDI RSC_TRK_W SDBM200W80_INV_BULK FN=2 WN=0.8U LN=0.03U 
+ MULTI=1 FP=4 WP=0.76U LP=0.03U
XINV6 Z8 VSSI VSSI VDDI VDDI CKPD SDBM200W80_INV_BULK FN=2 WN=0.76U LN=0.03U MULTI=1 
+ FP=2 WP=1.2U LP=0.03U
XINV5 CKP VSSI VSSI VDDI VDDI Z8 SDBM200W80_INV_BULK FN=1 WN=760N LN=0.03U MULTI=1 FP=1 
+ WP=1200N LP=0.03U
XI533 QLATCH VSSI VSSI VDDI VDDI NET096 SDBM200W80_INV_BULK FN=3 WN=0.87U LN=0.03U 
+ MULTI=1 FP=3 WP=1.2U LP=0.03U
XI635 TRKBL VSSI VSSI VDDI VDDI TRKBL_TM SDBM200W80_INV_BULK FN=1 WN=0.12U LN=30N 
+ MULTI=1 FP=1 WP=0.21U LP=30N
XI507 WLP_SAE VSSI VSSI VDDI VDDI NET0309 SDBM200W80_INV_BULK FN=1 WN=0.21U LN=0.03U 
+ MULTI=1 FP=1 WP=0.21U LP=0.03U
XI651 CKP_TRK VSSI VSSI VDDI VDDI NET0108 SDBM200W80_INV_BULK FN=2 WN=760N LN=0.03U 
+ MULTI=1 FP=2 WP=980N LP=0.03U
XI645 CKP_RED VSSI VSSI VDDI VDDI NET031 SDBM200W80_INV_BULK FN=1 WN=760N LN=0.03U 
+ MULTI=1 FP=1 WP=1200N LP=0.03U
XI647 NET031 VSSI VSSI VDDI VDDI CKPD_RED SDBM200W80_INV_BULK FN=4 WN=0.76U LN=0.03U 
+ MULTI=1 FP=4 WP=1.2U LP=0.03U
XI25 AXL VSSI VSSI VDDI VDDI D7 SDBM200W80_INV_BULK FN=1 WN=0.43U LN=0.03U MULTI=1 FP=2 
+ WP=0.32U LP=0.03U
XNAND3 CKP_TRK RTD_10 RTD_01_11 VSSI VSSI VDDI VDDI RTKB SDBM200W80_NAND3_BULK FN1=3 
+ WN1=1.2U LN1=30N FN2=3 WN2=1.2U LN2=30N FN3=3 WN3=1.2U LN3=30N FP3=2 
+ WP3=870N LP3=30N FP2=2 WP2=870N LP2=30N MULTI=1 FP1=2 WP1=870N LP1=30N
XTSEL_WT TRKBL1B VDDI VSSI NET0194 WV[0] WV[1] SDBM200W80_RESETD_TSEL_WT
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    COTH_M4_WOBIST_RED_DP_V3_H
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_COTH_M4_WOBIST_RED_DP_V3_H AWT AWT2 BLTRKWLDRV CKP CKP1 CKP2 CKPD 
+ CKPDCLK CKPD_RED CKP_RED CKP_TRK CLK QLATCH RSC RSC_TRK_H RSC_TRK_W RTSEL[0] 
+ RTSEL[1] TMA TMB TRKBL VDDI VHI VLO VSSI WEB2 WEB5B WLP_SAE WLP_SAEB 
+ WLP_SAE_TK WTSEL[0] WTSEL[1]
*.PININFO AWT:I CKP:I CKP1:I CKP2:I CKP_RED:I CKP_TRK:I CLK:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I TMA:I TMB:I WEB2:I WEB5B:I WTSEL[0]:I WTSEL[1]:I AWT2:O 
*.PININFO BLTRKWLDRV:O CKPD:O CKPDCLK:O CKPD_RED:O QLATCH:O RSC:O VHI:O VLO:O 
*.PININFO WLP_SAE:O WLP_SAEB:O RSC_TRK_H:B RSC_TRK_W:B TRKBL:B VDDI:B VSSI:B 
*.PININFO WLP_SAE_TK:B
XAWTD AWT AWT2 VDDI VSSI SDBM200W80_AWTD_M4
XRESETD BLTRKWLDRV CKP CKP1 CKP2 CKPD CKPDCLK CKPD_RED CKP_RED CKP_TRK CLK 
+ WLP_SAEB QLATCH RSC RSC_TRK_H RSC_TRK_W TMA TMB TRKBL VDDI VSSI WEB5B 
+ WLP_SAE WLP_SAE_TK RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] 
+ SDBM200W80_RESETD_M4_RED_DP_V3_H
XVHILO VDDI VHI VLO VSSI SDBM200W80_VHILO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CNT_CORE_M4_WOBIST_RED_DP_V3_H
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CNT_CORE_M4_WOBIST_RED_DP_V3_H AWT AWT2 BLTRKWLDRV CEB CK1B CK2 
+ CK2_TRK CKD CKP CKP2 CKP_RED CKP_TRK CLK DCLKA DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] QLATCH REDEN RSC RSC_TRK_H RSC_TRK_W RTSEL[0] RTSEL[1] TK 
+ TMA TMB TRKBL VDDI VHI VLO VSSI WEB WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] Y[0] Y[1]
*.PININFO AWT:I CEB:I CK1B:I CK2:I CK2_TRK:I CKP:I CKP2:I CKP_RED:I CKP_TRK:I 
*.PININFO CLK:I REDEN:I RTSEL[0]:I RTSEL[1]:I TMA:I TMB:I WEB:I WTSEL[0]:I 
*.PININFO WTSEL[1]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I Y[0]:I Y[1]:I AWT2:O BLTRKWLDRV:O CKD:O DCLKA:O 
*.PININFO DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O 
*.PININFO DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O 
*.PININFO DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O 
*.PININFO DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X3[0]:O DEC_X3[1]:O 
*.PININFO DEC_X3[2]:O DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O 
*.PININFO DEC_X3[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O 
*.PININFO DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O QLATCH:O RSC:O VHI:O VLO:O 
*.PININFO WLP_SAE:O WLP_SAEB:O RSC_TRK_H:B RSC_TRK_W:B TK:B TRKBL:B VDDI:B 
*.PININFO VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BLTRKWLDRV CKP CK2 CKP2 CKPD CKPDCLK CKPD_RED CKP_RED 
+ CKP_TRK CLK QLATCH RSC RSC_TRK_H RSC_TRK_W RTSEL[0] RTSEL[1] TMA TMB TRKBL 
+ VDDI VHI VLO VSSI WEB2 WEB5B WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ SDBM200W80_COTH_M4_WOBIST_RED_DP_V3_H
XCDEC CEB CK1B CK2 CK2_TRK CKD CKP CKPD CKPDCLK CKPD_RED CKP_RED DCLKA 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] REDEN VDDI VSSI WEB WEB2 WEB5B 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] Y[0] Y[1] 
+ SDBM200W80_CDEC_M4_WOBIST_RED_DP_V4
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CNT_WOBIST_M4_DP_0909_H
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CNT_WOBIST_M4_DP_0909_H AWT AWT2 BLTRKWLDRV CEBA CEBB CKD CLK DCLKA 
+ DCLK_L DCLK_R DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] DEC_X3[1] 
+ DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] 
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PHASESEL_L 
+ PHASESEL_R PTSEL[0] PTSEL[1] QCLKBA_L QCLKBA_R QCLKBB_L QCLKBB_R RSC_TRK_H 
+ RSC_TRK_W RTSEL[0] RTSEL[1] TMA TMB TRKBL VDDI VHI VLO VSSI WEBA WEBB 
+ WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] XA[9] XA[8] XA[7] XA[6] XA[5] 
+ XA[4] XA[3] XA[2] XA[1] XA[0] XB[9] XB[8] XB[7] XB[6] XB[5] XB[4] XB[3] 
+ XB[2] XB[1] XB[0] YA[1] YA[0] YB[1] YB[0]
*.PININFO AWT:I CEBA:I CEBB:I CLK:I PTSEL[0]:I PTSEL[1]:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I TMA:I TMB:I WEBA:I WEBB:I WLP_SAE_TK:I WTSEL[0]:I 
*.PININFO WTSEL[1]:I XA[9]:I XA[8]:I XA[7]:I XA[6]:I XA[5]:I XA[4]:I XA[3]:I 
*.PININFO XA[2]:I XA[1]:I XA[0]:I XB[9]:I XB[8]:I XB[7]:I XB[6]:I XB[5]:I 
*.PININFO XB[4]:I XB[3]:I XB[2]:I XB[1]:I XB[0]:I YA[1]:I YA[0]:I YB[1]:I 
*.PININFO YB[0]:I AWT2:O BLTRKWLDRV:O CKD:O DCLKA:O DCLK_L:O DCLK_R:O 
*.PININFO DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O 
*.PININFO DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O 
*.PININFO DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O 
*.PININFO DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X3[0]:O DEC_X3[1]:O 
*.PININFO DEC_X3[2]:O DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O 
*.PININFO DEC_X3[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O 
*.PININFO DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PHASESEL_L:O PHASESEL_R:O 
*.PININFO QCLKBA_L:O QCLKBA_R:O QCLKBB_L:O QCLKBB_R:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O RSC_TRK_H:B RSC_TRK_W:B TRKBL:B VDDI:B VSSI:B
XCNT_WRAPPER YA[1] YA[0] XA[9] XA[8] XA[7] XA[6] XA[5] XA[4] XA[3] XA[2] XA[1] 
+ XA[0] YB[1] YB[0] XB[9] XB[8] XB[7] XB[6] XB[5] XB[4] XB[3] XB[2] XB[1] 
+ XB[0] X[9] X[8] X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] Y[1] Y[0] CEBA CEBB 
+ CEB CKP1 CKP1_TRK CKP2 CKPB1 CKP_EN CKP_RSTB CKP_TRK CKT CLK CKP CKP_RED 
+ DCLK_L DCLK_R QLATCH PHASESEL_L PHASESEL_R PTSEL[0] PTSEL[1] QCLKBA_L 
+ QCLKBA_R QCLKBB_L QCLKBB_R VLO VHI VDDI VSSI WEBA WEBB WEB SDBM200W80_CNT_WP_M4_V5
XI27 CKP1 VSSI VSSI VDDI VDDI CK1B SDBM200W80_INV_BULK FN=3 WN=0.65U LN=0.03U MULTI=1 
+ FP=3 WP=0.76U LP=0.03U
XCNT_CORE AWT AWT2 BLTRKWLDRV CEB CK1B CKP1 CKP1_TRK CKD CKP CKP2 CKP_RED 
+ CKP_TRK CLK DCLKA DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ QLATCH VLO CKP_RSTB RSC_TRK_H RSC_TRK_W RTSEL[0] RTSEL[1] NET23 TMA TMB 
+ TRKBL VDDI VHI VLO VSSI WEB WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] Y[0] Y[1] 
+ SDBM200W80_CNT_CORE_M4_WOBIST_RED_DP_V3_H
.ENDS

************************************************************************
* LIBRARY NAME: N28HPM_DP_LEAFCELLS
* CELL NAME:    CNT_WOBIST_M4_DP_IOX10_HALF
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT SDBM200W80_CNT_WOBIST_M4_DP_IOX10_HALF AWT AWT2 BLTRKWLDRV BWEBA[0] BWEBA[1] 
+ BWEBA[2] BWEBA[3] BWEBA[4] BWEBA[5] BWEBA[6] BWEBA[7] BWEBA_L BWEBA_R 
+ BWEBB[0] BWEBB[1] BWEBB[2] BWEBB[3] BWEBB[4] BWEBB[5] BWEBB[6] BWEBB[7] 
+ BWEBB_L BWEBB_R CEBA CEBB CKD CLK DA[0] DA[1] DA[2] DA[3] DA[4] DA[5] DA[6] 
+ DA[7] DA_L DA_R DB[0] DB[1] DB[2] DB[3] DB[4] DB[5] DB[6] DB[7] DB_L DB_R 
+ DCLKA DCLK_L DCLK_R DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBLB[0] GBLB[1] 
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB_L GBLB_R GBL_L GBL_R 
+ GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GWB[0] GWB[1] GWB[2] GWB[3] 
+ GWB[4] GWB[5] GWB[6] GWB[7] GWB_L GWB_R GW_L GW_R PHASESEL_L PHASESEL_R 
+ PTSEL[0] PTSEL[1] QA[0] QA[1] QA[2] QA[3] QA[4] QA[5] QA[6] QA[7] QA_L QA_R 
+ QB[0] QB[1] QB[2] QB[3] QB[4] QB[5] QB[6] QB[7] QB_L QB_R QLATCH_AB_L 
+ QLATCH_AB_R QLATCH_BB_L QLATCH_BB_R RSC_TRK_H RSC_TRK_W RTSEL[0] RTSEL[1] 
+ TMA TMB TRKBL VDDI VHI VLO VSSI WEBA WEBB WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] XA[0] XA[1] XA[2] XA[3] XA[4] XA[5] XA[6] XA[7] XA[8] 
+ XA[9] XB[0] XB[1] XB[2] XB[3] XB[4] XB[5] XB[6] XB[7] XB[8] XB[9] YA[0] 
+ YA[1] YB[0] YB[1]
*.PININFO AWT:I BWEBA[0]:I BWEBA[1]:I BWEBA[2]:I BWEBA[3]:I BWEBA[4]:I 
*.PININFO BWEBA[5]:I BWEBA[6]:I BWEBA[7]:I BWEBA_L:I BWEBA_R:I BWEBB[0]:I 
*.PININFO BWEBB[1]:I BWEBB[2]:I BWEBB[3]:I BWEBB[4]:I BWEBB[5]:I BWEBB[6]:I 
*.PININFO BWEBB[7]:I BWEBB_L:I BWEBB_R:I CEBA:I CEBB:I CLK:I DA[0]:I DA[1]:I 
*.PININFO DA[2]:I DA[3]:I DA[4]:I DA[5]:I DA[6]:I DA[7]:I DA_L:I DA_R:I 
*.PININFO DB[0]:I DB[1]:I DB[2]:I DB[3]:I DB[4]:I DB[5]:I DB[6]:I DB[7]:I 
*.PININFO DB_L:I DB_R:I PTSEL[0]:I PTSEL[1]:I RTSEL[0]:I RTSEL[1]:I TMA:I 
*.PININFO TMB:I WEBA:I WEBB:I WTSEL[0]:I WTSEL[1]:I XA[0]:I XA[1]:I XA[2]:I 
*.PININFO XA[3]:I XA[4]:I XA[5]:I XA[6]:I XA[7]:I XA[8]:I XA[9]:I XB[0]:I 
*.PININFO XB[1]:I XB[2]:I XB[3]:I XB[4]:I XB[5]:I XB[6]:I XB[7]:I XB[8]:I 
*.PININFO XB[9]:I YA[0]:I YA[1]:I YB[0]:I YB[1]:I QA[0]:O QA[1]:O QA[2]:O 
*.PININFO QA[3]:O QA[4]:O QA[5]:O QA[6]:O QA[7]:O QA_L:O QA_R:O QB[0]:O 
*.PININFO QB[1]:O QB[2]:O QB[3]:O QB[4]:O QB[5]:O QB[6]:O QB[7]:O QB_L:O 
*.PININFO QB_R:O AWT2:B BLTRKWLDRV:B CKD:B DCLKA:B DCLK_L:B DCLK_R:B 
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X3[0]:B DEC_X3[1]:B 
*.PININFO DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B 
*.PININFO DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B 
*.PININFO DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B 
*.PININFO GBL[4]:B GBL[5]:B GBL[6]:B GBL[7]:B GBLB[0]:B GBLB[1]:B GBLB[2]:B 
*.PININFO GBLB[3]:B GBLB[4]:B GBLB[5]:B GBLB[6]:B GBLB[7]:B GBLB_L:B GBLB_R:B 
*.PININFO GBL_L:B GBL_R:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B GW[4]:B GW[5]:B 
*.PININFO GW[6]:B GW[7]:B GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B GWB[4]:B 
*.PININFO GWB[5]:B GWB[6]:B GWB[7]:B GWB_L:B GWB_R:B GW_L:B GW_R:B 
*.PININFO PHASESEL_L:B PHASESEL_R:B QLATCH_AB_L:B QLATCH_AB_R:B QLATCH_BB_L:B 
*.PININFO QLATCH_BB_R:B RSC_TRK_H:B RSC_TRK_W:B TRKBL:B VDDI:B VHI:B VLO:B 
*.PININFO VSSI:B WLP_SAE:B WLP_SAEB:B WLP_SAE_TK:B
XMIO[5] AWT2 BWEBA_R BWEBB_R CKD DA_R DB_R DCLK_R DCLKA GBL_R GBLB_R GW_R 
+ GWB_R PHASESEL_R QA_R QB_R QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI 
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[6] AWT2 BWEBA[4] BWEBB[4] CKD DA[4] DB[4] DCLK_R DCLKA GBL[4] GBLB[4] 
+ GW[4] GWB[4] PHASESEL_R QA[4] QB[4] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI 
+ VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[7] AWT2 BWEBA[5] BWEBB[5] CKD DA[5] DB[5] DCLK_R DCLKA GBL[5] GBLB[5] 
+ GW[5] GWB[5] PHASESEL_R QA[5] QB[5] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI 
+ VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[8] AWT2 BWEBA[6] BWEBB[6] CKD DA[6] DB[6] DCLK_R DCLKA GBL[6] GBLB[6] 
+ GW[6] GWB[6] PHASESEL_R QA[6] QB[6] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI 
+ VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[9] AWT2 BWEBA[7] BWEBB[7] CKD DA[7] DB[7] DCLK_R DCLKA GBL[7] GBLB[7] 
+ GW[7] GWB[7] PHASESEL_R QA[7] QB[7] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI 
+ VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[0] AWT2 BWEBA[0] BWEBB[0] CKD DA[0] DB[0] DCLK_L DCLKA GBL[0] GBLB[0] 
+ GW[0] GWB[0] PHASESEL_L QA[0] QB[0] QLATCH_AB_L QLATCH_BB_L NET017 VDDI VSSI 
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[1] AWT2 BWEBA[1] BWEBB[1] CKD DA[1] DB[1] DCLK_L DCLKA GBL[1] GBLB[1] 
+ GW[1] GWB[1] PHASESEL_L QA[1] QB[1] QLATCH_AB_L QLATCH_BB_L NET017 VDDI VSSI 
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[2] AWT2 BWEBA[2] BWEBB[2] CKD DA[2] DB[2] DCLK_L DCLKA GBL[2] GBLB[2] 
+ GW[2] GWB[2] PHASESEL_L QA[2] QB[2] QLATCH_AB_L QLATCH_BB_L NET017 VDDI VSSI 
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[3] AWT2 BWEBA[3] BWEBB[3] CKD DA[3] DB[3] DCLK_L DCLKA GBL[3] GBLB[3] 
+ GW[3] GWB[3] PHASESEL_L QA[3] QB[3] QLATCH_AB_L QLATCH_BB_L NET017 VDDI VSSI 
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XMIO[4] AWT2 BWEBA_L BWEBB_L CKD DA_L DB_L DCLK_L DCLKA GBL_L GBLB_L GW_L 
+ GWB_L PHASESEL_L QA_L QB_L QLATCH_AB_L QLATCH_BB_L NET017 VDDI VSSI WLP_SAEB 
+ SDBM200W80_IO_WOBIST_DP
XCNT AWT AWT2 BLTRKWLDRV CEBA CEBB CKD CLK DCLKA DCLK_L DCLK_R DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PHASESEL_L PHASESEL_R PTSEL[0] PTSEL[1] 
+ QLATCH_AB_L QLATCH_AB_R QLATCH_BB_L QLATCH_BB_R RSC_TRK_H RSC_TRK_W RTSEL[0] 
+ RTSEL[1] TMA TMB TRKBL VDDI VHI VLO VSSI WEBA WEBB WLP_SAE WLP_SAEB 
+ WLP_SAE_TK WTSEL[0] WTSEL[1] XA[9] XA[8] XA[7] XA[6] XA[5] XA[4] XA[3] XA[2] 
+ XA[1] XA[0] XB[9] XB[8] XB[7] XB[6] XB[5] XB[4] XB[3] XB[2] XB[1] XB[0] 
+ YA[1] YA[0] YB[1] YB[0] SDBM200W80_CNT_WOBIST_M4_DP_0909_H
.ENDS




**** End of leaf cells

.SUBCKT SDBM200W80_CELL_ARR_X BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7]
+ BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18]
+ BL[19] BL[20] BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29]
+ BL[30] BL[31] BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40]
+ BL[41] BL[42] BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51]
+ BL[52] BL[53] BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62]
+ BL[63] BL[64] BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73]
+ BL[74] BL[75] BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84]
+ BL[85] BL[86] BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95]
+ BL[96] BL[97] BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105]
+ BL[106] BL[107] BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114]
+ BL[115] BL[116] BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123]
+ BL[124] BL[125] BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132]
+ BL[133] BL[134] BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141]
+ BL[142] BL[143] BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150]
+ BL[151] BL[152] BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159]
+ BL[160] BL[161] BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168]
+ BL[169] BL[170] BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177]
+ BL[178] BL[179] BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186]
+ BL[187] BL[188] BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195]
+ BL[196] BL[197] BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204]
+ BL[205] BL[206] BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213]
+ BL[214] BL[215] BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222]
+ BL[223] BL[224] BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231]
+ BL[232] BL[233] BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240]
+ BL[241] BL[242] BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249]
+ BL[250] BL[251] BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258]
+ BL[259] BL[260] BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267]
+ BL[268] BL[269] BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276]
+ BL[277] BL[278] BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285]
+ BL[286] BL[287] BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294]
+ BL[295] BL[296] BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303]
+ BL[304] BL[305] BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312]
+ BL[313] BL[314] BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321]
+ BL[322] BL[323] BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330]
+ BL[331] BL[332] BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339]
+ BL[340] BL[341] BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348]
+ BL[349] BL[350] BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357]
+ BL[358] BL[359] BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366]
+ BL[367] BL[368] BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375]
+ BL[376] BL[377] BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384]
+ BL[385] BL[386] BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393]
+ BL[394] BL[395] BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402]
+ BL[403] BL[404] BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411]
+ BL[412] BL[413] BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420]
+ BL[421] BL[422] BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429]
+ BL[430] BL[431] BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438]
+ BL[439] BL[440] BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447]
+ BL[448] BL[449] BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456]
+ BL[457] BL[458] BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465]
+ BL[466] BL[467] BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474]
+ BL[475] BL[476] BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483]
+ BL[484] BL[485] BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492]
+ BL[493] BL[494] BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501]
+ BL[502] BL[503] BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510]
+ BL[511] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9]
+ BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18]
+ BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27]
+ BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36]
+ BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45]
+ BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54]
+ BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63]
+ BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72]
+ BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81]
+ BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90]
+ BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99]
+ BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107]
+ BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115]
+ BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123]
+ BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131]
+ BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139]
+ BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147]
+ BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155]
+ BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163]
+ BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171]
+ BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179]
+ BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187]
+ BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195]
+ BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203]
+ BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211]
+ BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219]
+ BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227]
+ BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235]
+ BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243]
+ BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251]
+ BLB[252] BLB[253] BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259]
+ BLB[260] BLB[261] BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267]
+ BLB[268] BLB[269] BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275]
+ BLB[276] BLB[277] BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283]
+ BLB[284] BLB[285] BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291]
+ BLB[292] BLB[293] BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299]
+ BLB[300] BLB[301] BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307]
+ BLB[308] BLB[309] BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315]
+ BLB[316] BLB[317] BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323]
+ BLB[324] BLB[325] BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331]
+ BLB[332] BLB[333] BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339]
+ BLB[340] BLB[341] BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347]
+ BLB[348] BLB[349] BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355]
+ BLB[356] BLB[357] BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363]
+ BLB[364] BLB[365] BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371]
+ BLB[372] BLB[373] BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379]
+ BLB[380] BLB[381] BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387]
+ BLB[388] BLB[389] BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395]
+ BLB[396] BLB[397] BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403]
+ BLB[404] BLB[405] BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411]
+ BLB[412] BLB[413] BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419]
+ BLB[420] BLB[421] BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427]
+ BLB[428] BLB[429] BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435]
+ BLB[436] BLB[437] BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443]
+ BLB[444] BLB[445] BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451]
+ BLB[452] BLB[453] BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459]
+ BLB[460] BLB[461] BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467]
+ BLB[468] BLB[469] BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475]
+ BLB[476] BLB[477] BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483]
+ BLB[484] BLB[485] BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491]
+ BLB[492] BLB[493] BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499]
+ BLB[500] BLB[501] BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507]
+ BLB[508] BLB[509] BLB[510] BLB[511] WL[0] WL[1] VDDI VSSI GBL[0] GBL[1] GBL[2]
+ GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12]
+ GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21]
+ GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30]
+ GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39]
+ GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48]
+ GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57]
+ GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66]
+ GBL[67] GBL[68] GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75]
+ GBL[76] GBL[77] GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84]
+ GBL[85] GBL[86] GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93]
+ GBL[94] GBL[95] GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102]
+ GBL[103] GBL[104] GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110]
+ GBL[111] GBL[112] GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118]
+ GBL[119] GBL[120] GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126]
+ GBL[127] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7]
+ GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16]
+ GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24]
+ GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32]
+ GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40]
+ GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48]
+ GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56]
+ GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64]
+ GBLB[65] GBLB[66] GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72]
+ GBLB[73] GBLB[74] GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80]
+ GBLB[81] GBLB[82] GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88]
+ GBLB[89] GBLB[90] GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96]
+ GBLB[97] GBLB[98] GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104]
+ GBLB[105] GBLB[106] GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111]
+ GBLB[112] GBLB[113] GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118]
+ GBLB[119] GBLB[120] GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125]
+ GBLB[126] GBLB[127] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8]
+ GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19]
+ GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30]
+ GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41]
+ GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52]
+ GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63]
+ GW[64] GW[65] GW[66] GW[67] GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74]
+ GW[75] GW[76] GW[77] GW[78] GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85]
+ GW[86] GW[87] GW[88] GW[89] GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96]
+ GW[97] GW[98] GW[99] GW[100] GW[101] GW[102] GW[103] GW[104] GW[105] GW[106]
+ GW[107] GW[108] GW[109] GW[110] GW[111] GW[112] GW[113] GW[114] GW[115]
+ GW[116] GW[117] GW[118] GW[119] GW[120] GW[121] GW[122] GW[123] GW[124]
+ GW[125] GW[126] GW[127] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] GWB[64] GWB[65] GWB[66] GWB[67] GWB[68] GWB[69] GWB[70]
+ GWB[71] GWB[72] GWB[73] GWB[74] GWB[75] GWB[76] GWB[77] GWB[78] GWB[79]
+ GWB[80] GWB[81] GWB[82] GWB[83] GWB[84] GWB[85] GWB[86] GWB[87] GWB[88]
+ GWB[89] GWB[90] GWB[91] GWB[92] GWB[93] GWB[94] GWB[95] GWB[96] GWB[97]
+ GWB[98] GWB[99] GWB[100] GWB[101] GWB[102] GWB[103] GWB[104] GWB[105] GWB[106]
+ GWB[107] GWB[108] GWB[109] GWB[110] GWB[111] GWB[112] GWB[113] GWB[114]
+ GWB[115] GWB[116] GWB[117] GWB[118] GWB[119] GWB[120] GWB[121] GWB[122]
+ GWB[123] GWB[124] GWB[125] GWB[126] GWB[127]
XMCB_0 BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL[0] GBLB[0] GW[0]
+ GWB[0] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_1 BL[4] BL[5] BL[6] BL[7] BLB[4] BLB[5] BLB[6] BLB[7] GBL[1] GBLB[1] GW[1]
+ GWB[1] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_2 BL[8] BL[9] BL[10] BL[11] BLB[8] BLB[9] BLB[10] BLB[11] GBL[2] GBLB[2]
+ GW[2] GWB[2] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_3 BL[12] BL[13] BL[14] BL[15] BLB[12] BLB[13] BLB[14] BLB[15] GBL[3]
+ GBLB[3] GW[3] GWB[3] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_4 BL[16] BL[17] BL[18] BL[19] BLB[16] BLB[17] BLB[18] BLB[19] GBL[4]
+ GBLB[4] GW[4] GWB[4] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_5 BL[20] BL[21] BL[22] BL[23] BLB[20] BLB[21] BLB[22] BLB[23] GBL[5]
+ GBLB[5] GW[5] GWB[5] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_6 BL[24] BL[25] BL[26] BL[27] BLB[24] BLB[25] BLB[26] BLB[27] GBL[6]
+ GBLB[6] GW[6] GWB[6] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_7 BL[28] BL[29] BL[30] BL[31] BLB[28] BLB[29] BLB[30] BLB[31] GBL[7]
+ GBLB[7] GW[7] GWB[7] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_8 BL[32] BL[33] BL[34] BL[35] BLB[32] BLB[33] BLB[34] BLB[35] GBL[8]
+ GBLB[8] GW[8] GWB[8] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_9 BL[36] BL[37] BL[38] BL[39] BLB[36] BLB[37] BLB[38] BLB[39] GBL[9]
+ GBLB[9] GW[9] GWB[9] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_10 BL[40] BL[41] BL[42] BL[43] BLB[40] BLB[41] BLB[42] BLB[43] GBL[10]
+ GBLB[10] GW[10] GWB[10] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_11 BL[44] BL[45] BL[46] BL[47] BLB[44] BLB[45] BLB[46] BLB[47] GBL[11]
+ GBLB[11] GW[11] GWB[11] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_12 BL[48] BL[49] BL[50] BL[51] BLB[48] BLB[49] BLB[50] BLB[51] GBL[12]
+ GBLB[12] GW[12] GWB[12] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_13 BL[52] BL[53] BL[54] BL[55] BLB[52] BLB[53] BLB[54] BLB[55] GBL[13]
+ GBLB[13] GW[13] GWB[13] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_14 BL[56] BL[57] BL[58] BL[59] BLB[56] BLB[57] BLB[58] BLB[59] GBL[14]
+ GBLB[14] GW[14] GWB[14] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_15 BL[60] BL[61] BL[62] BL[63] BLB[60] BLB[61] BLB[62] BLB[63] GBL[15]
+ GBLB[15] GW[15] GWB[15] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_16 BL[64] BL[65] BL[66] BL[67] BLB[64] BLB[65] BLB[66] BLB[67] GBL[16]
+ GBLB[16] GW[16] GWB[16] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_17 BL[68] BL[69] BL[70] BL[71] BLB[68] BLB[69] BLB[70] BLB[71] GBL[17]
+ GBLB[17] GW[17] GWB[17] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_18 BL[72] BL[73] BL[74] BL[75] BLB[72] BLB[73] BLB[74] BLB[75] GBL[18]
+ GBLB[18] GW[18] GWB[18] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_19 BL[76] BL[77] BL[78] BL[79] BLB[76] BLB[77] BLB[78] BLB[79] GBL[19]
+ GBLB[19] GW[19] GWB[19] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_20 BL[80] BL[81] BL[82] BL[83] BLB[80] BLB[81] BLB[82] BLB[83] GBL[20]
+ GBLB[20] GW[20] GWB[20] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_21 BL[84] BL[85] BL[86] BL[87] BLB[84] BLB[85] BLB[86] BLB[87] GBL[21]
+ GBLB[21] GW[21] GWB[21] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_22 BL[88] BL[89] BL[90] BL[91] BLB[88] BLB[89] BLB[90] BLB[91] GBL[22]
+ GBLB[22] GW[22] GWB[22] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_23 BL[92] BL[93] BL[94] BL[95] BLB[92] BLB[93] BLB[94] BLB[95] GBL[23]
+ GBLB[23] GW[23] GWB[23] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_24 BL[96] BL[97] BL[98] BL[99] BLB[96] BLB[97] BLB[98] BLB[99] GBL[24]
+ GBLB[24] GW[24] GWB[24] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_25 BL[100] BL[101] BL[102] BL[103] BLB[100] BLB[101] BLB[102] BLB[103]
+ GBL[25] GBLB[25] GW[25] GWB[25] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_26 BL[104] BL[105] BL[106] BL[107] BLB[104] BLB[105] BLB[106] BLB[107]
+ GBL[26] GBLB[26] GW[26] GWB[26] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_27 BL[108] BL[109] BL[110] BL[111] BLB[108] BLB[109] BLB[110] BLB[111]
+ GBL[27] GBLB[27] GW[27] GWB[27] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_28 BL[112] BL[113] BL[114] BL[115] BLB[112] BLB[113] BLB[114] BLB[115]
+ GBL[28] GBLB[28] GW[28] GWB[28] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_29 BL[116] BL[117] BL[118] BL[119] BLB[116] BLB[117] BLB[118] BLB[119]
+ GBL[29] GBLB[29] GW[29] GWB[29] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_30 BL[120] BL[121] BL[122] BL[123] BLB[120] BLB[121] BLB[122] BLB[123]
+ GBL[30] GBLB[30] GW[30] GWB[30] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_31 BL[124] BL[125] BL[126] BL[127] BLB[124] BLB[125] BLB[126] BLB[127]
+ GBL[31] GBLB[31] GW[31] GWB[31] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_32 BL[128] BL[129] BL[130] BL[131] BLB[128] BLB[129] BLB[130] BLB[131]
+ GBL[32] GBLB[32] GW[32] GWB[32] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_33 BL[132] BL[133] BL[134] BL[135] BLB[132] BLB[133] BLB[134] BLB[135]
+ GBL[33] GBLB[33] GW[33] GWB[33] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_34 BL[136] BL[137] BL[138] BL[139] BLB[136] BLB[137] BLB[138] BLB[139]
+ GBL[34] GBLB[34] GW[34] GWB[34] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_35 BL[140] BL[141] BL[142] BL[143] BLB[140] BLB[141] BLB[142] BLB[143]
+ GBL[35] GBLB[35] GW[35] GWB[35] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_36 BL[144] BL[145] BL[146] BL[147] BLB[144] BLB[145] BLB[146] BLB[147]
+ GBL[36] GBLB[36] GW[36] GWB[36] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_37 BL[148] BL[149] BL[150] BL[151] BLB[148] BLB[149] BLB[150] BLB[151]
+ GBL[37] GBLB[37] GW[37] GWB[37] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_38 BL[152] BL[153] BL[154] BL[155] BLB[152] BLB[153] BLB[154] BLB[155]
+ GBL[38] GBLB[38] GW[38] GWB[38] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_39 BL[156] BL[157] BL[158] BL[159] BLB[156] BLB[157] BLB[158] BLB[159]
+ GBL[39] GBLB[39] GW[39] GWB[39] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_40 BL[160] BL[161] BL[162] BL[163] BLB[160] BLB[161] BLB[162] BLB[163]
+ GBL[40] GBLB[40] GW[40] GWB[40] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_41 BL[164] BL[165] BL[166] BL[167] BLB[164] BLB[165] BLB[166] BLB[167]
+ GBL[41] GBLB[41] GW[41] GWB[41] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_42 BL[168] BL[169] BL[170] BL[171] BLB[168] BLB[169] BLB[170] BLB[171]
+ GBL[42] GBLB[42] GW[42] GWB[42] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_43 BL[172] BL[173] BL[174] BL[175] BLB[172] BLB[173] BLB[174] BLB[175]
+ GBL[43] GBLB[43] GW[43] GWB[43] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_44 BL[176] BL[177] BL[178] BL[179] BLB[176] BLB[177] BLB[178] BLB[179]
+ GBL[44] GBLB[44] GW[44] GWB[44] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_45 BL[180] BL[181] BL[182] BL[183] BLB[180] BLB[181] BLB[182] BLB[183]
+ GBL[45] GBLB[45] GW[45] GWB[45] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_46 BL[184] BL[185] BL[186] BL[187] BLB[184] BLB[185] BLB[186] BLB[187]
+ GBL[46] GBLB[46] GW[46] GWB[46] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_47 BL[188] BL[189] BL[190] BL[191] BLB[188] BLB[189] BLB[190] BLB[191]
+ GBL[47] GBLB[47] GW[47] GWB[47] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_48 BL[192] BL[193] BL[194] BL[195] BLB[192] BLB[193] BLB[194] BLB[195]
+ GBL[48] GBLB[48] GW[48] GWB[48] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_49 BL[196] BL[197] BL[198] BL[199] BLB[196] BLB[197] BLB[198] BLB[199]
+ GBL[49] GBLB[49] GW[49] GWB[49] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_50 BL[200] BL[201] BL[202] BL[203] BLB[200] BLB[201] BLB[202] BLB[203]
+ GBL[50] GBLB[50] GW[50] GWB[50] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_51 BL[204] BL[205] BL[206] BL[207] BLB[204] BLB[205] BLB[206] BLB[207]
+ GBL[51] GBLB[51] GW[51] GWB[51] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_52 BL[208] BL[209] BL[210] BL[211] BLB[208] BLB[209] BLB[210] BLB[211]
+ GBL[52] GBLB[52] GW[52] GWB[52] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_53 BL[212] BL[213] BL[214] BL[215] BLB[212] BLB[213] BLB[214] BLB[215]
+ GBL[53] GBLB[53] GW[53] GWB[53] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_54 BL[216] BL[217] BL[218] BL[219] BLB[216] BLB[217] BLB[218] BLB[219]
+ GBL[54] GBLB[54] GW[54] GWB[54] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_55 BL[220] BL[221] BL[222] BL[223] BLB[220] BLB[221] BLB[222] BLB[223]
+ GBL[55] GBLB[55] GW[55] GWB[55] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_56 BL[224] BL[225] BL[226] BL[227] BLB[224] BLB[225] BLB[226] BLB[227]
+ GBL[56] GBLB[56] GW[56] GWB[56] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_57 BL[228] BL[229] BL[230] BL[231] BLB[228] BLB[229] BLB[230] BLB[231]
+ GBL[57] GBLB[57] GW[57] GWB[57] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_58 BL[232] BL[233] BL[234] BL[235] BLB[232] BLB[233] BLB[234] BLB[235]
+ GBL[58] GBLB[58] GW[58] GWB[58] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_59 BL[236] BL[237] BL[238] BL[239] BLB[236] BLB[237] BLB[238] BLB[239]
+ GBL[59] GBLB[59] GW[59] GWB[59] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_60 BL[240] BL[241] BL[242] BL[243] BLB[240] BLB[241] BLB[242] BLB[243]
+ GBL[60] GBLB[60] GW[60] GWB[60] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_61 BL[244] BL[245] BL[246] BL[247] BLB[244] BLB[245] BLB[246] BLB[247]
+ GBL[61] GBLB[61] GW[61] GWB[61] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_62 BL[248] BL[249] BL[250] BL[251] BLB[248] BLB[249] BLB[250] BLB[251]
+ GBL[62] GBLB[62] GW[62] GWB[62] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_63 BL[252] BL[253] BL[254] BL[255] BLB[252] BLB[253] BLB[254] BLB[255]
+ GBL[63] GBLB[63] GW[63] GWB[63] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_64 BL[256] BL[257] BL[258] BL[259] BLB[256] BLB[257] BLB[258] BLB[259]
+ GBL[64] GBLB[64] GW[64] GWB[64] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_65 BL[260] BL[261] BL[262] BL[263] BLB[260] BLB[261] BLB[262] BLB[263]
+ GBL[65] GBLB[65] GW[65] GWB[65] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_66 BL[264] BL[265] BL[266] BL[267] BLB[264] BLB[265] BLB[266] BLB[267]
+ GBL[66] GBLB[66] GW[66] GWB[66] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_67 BL[268] BL[269] BL[270] BL[271] BLB[268] BLB[269] BLB[270] BLB[271]
+ GBL[67] GBLB[67] GW[67] GWB[67] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_68 BL[272] BL[273] BL[274] BL[275] BLB[272] BLB[273] BLB[274] BLB[275]
+ GBL[68] GBLB[68] GW[68] GWB[68] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_69 BL[276] BL[277] BL[278] BL[279] BLB[276] BLB[277] BLB[278] BLB[279]
+ GBL[69] GBLB[69] GW[69] GWB[69] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_70 BL[280] BL[281] BL[282] BL[283] BLB[280] BLB[281] BLB[282] BLB[283]
+ GBL[70] GBLB[70] GW[70] GWB[70] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_71 BL[284] BL[285] BL[286] BL[287] BLB[284] BLB[285] BLB[286] BLB[287]
+ GBL[71] GBLB[71] GW[71] GWB[71] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_72 BL[288] BL[289] BL[290] BL[291] BLB[288] BLB[289] BLB[290] BLB[291]
+ GBL[72] GBLB[72] GW[72] GWB[72] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_73 BL[292] BL[293] BL[294] BL[295] BLB[292] BLB[293] BLB[294] BLB[295]
+ GBL[73] GBLB[73] GW[73] GWB[73] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_74 BL[296] BL[297] BL[298] BL[299] BLB[296] BLB[297] BLB[298] BLB[299]
+ GBL[74] GBLB[74] GW[74] GWB[74] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_75 BL[300] BL[301] BL[302] BL[303] BLB[300] BLB[301] BLB[302] BLB[303]
+ GBL[75] GBLB[75] GW[75] GWB[75] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_76 BL[304] BL[305] BL[306] BL[307] BLB[304] BLB[305] BLB[306] BLB[307]
+ GBL[76] GBLB[76] GW[76] GWB[76] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_77 BL[308] BL[309] BL[310] BL[311] BLB[308] BLB[309] BLB[310] BLB[311]
+ GBL[77] GBLB[77] GW[77] GWB[77] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_78 BL[312] BL[313] BL[314] BL[315] BLB[312] BLB[313] BLB[314] BLB[315]
+ GBL[78] GBLB[78] GW[78] GWB[78] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_79 BL[316] BL[317] BL[318] BL[319] BLB[316] BLB[317] BLB[318] BLB[319]
+ GBL[79] GBLB[79] GW[79] GWB[79] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_80 BL[320] BL[321] BL[322] BL[323] BLB[320] BLB[321] BLB[322] BLB[323]
+ GBL[80] GBLB[80] GW[80] GWB[80] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_81 BL[324] BL[325] BL[326] BL[327] BLB[324] BLB[325] BLB[326] BLB[327]
+ GBL[81] GBLB[81] GW[81] GWB[81] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_82 BL[328] BL[329] BL[330] BL[331] BLB[328] BLB[329] BLB[330] BLB[331]
+ GBL[82] GBLB[82] GW[82] GWB[82] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_83 BL[332] BL[333] BL[334] BL[335] BLB[332] BLB[333] BLB[334] BLB[335]
+ GBL[83] GBLB[83] GW[83] GWB[83] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_84 BL[336] BL[337] BL[338] BL[339] BLB[336] BLB[337] BLB[338] BLB[339]
+ GBL[84] GBLB[84] GW[84] GWB[84] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_85 BL[340] BL[341] BL[342] BL[343] BLB[340] BLB[341] BLB[342] BLB[343]
+ GBL[85] GBLB[85] GW[85] GWB[85] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_86 BL[344] BL[345] BL[346] BL[347] BLB[344] BLB[345] BLB[346] BLB[347]
+ GBL[86] GBLB[86] GW[86] GWB[86] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_87 BL[348] BL[349] BL[350] BL[351] BLB[348] BLB[349] BLB[350] BLB[351]
+ GBL[87] GBLB[87] GW[87] GWB[87] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_88 BL[352] BL[353] BL[354] BL[355] BLB[352] BLB[353] BLB[354] BLB[355]
+ GBL[88] GBLB[88] GW[88] GWB[88] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_89 BL[356] BL[357] BL[358] BL[359] BLB[356] BLB[357] BLB[358] BLB[359]
+ GBL[89] GBLB[89] GW[89] GWB[89] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_90 BL[360] BL[361] BL[362] BL[363] BLB[360] BLB[361] BLB[362] BLB[363]
+ GBL[90] GBLB[90] GW[90] GWB[90] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_91 BL[364] BL[365] BL[366] BL[367] BLB[364] BLB[365] BLB[366] BLB[367]
+ GBL[91] GBLB[91] GW[91] GWB[91] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_92 BL[368] BL[369] BL[370] BL[371] BLB[368] BLB[369] BLB[370] BLB[371]
+ GBL[92] GBLB[92] GW[92] GWB[92] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_93 BL[372] BL[373] BL[374] BL[375] BLB[372] BLB[373] BLB[374] BLB[375]
+ GBL[93] GBLB[93] GW[93] GWB[93] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_94 BL[376] BL[377] BL[378] BL[379] BLB[376] BLB[377] BLB[378] BLB[379]
+ GBL[94] GBLB[94] GW[94] GWB[94] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_95 BL[380] BL[381] BL[382] BL[383] BLB[380] BLB[381] BLB[382] BLB[383]
+ GBL[95] GBLB[95] GW[95] GWB[95] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_96 BL[384] BL[385] BL[386] BL[387] BLB[384] BLB[385] BLB[386] BLB[387]
+ GBL[96] GBLB[96] GW[96] GWB[96] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_97 BL[388] BL[389] BL[390] BL[391] BLB[388] BLB[389] BLB[390] BLB[391]
+ GBL[97] GBLB[97] GW[97] GWB[97] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_98 BL[392] BL[393] BL[394] BL[395] BLB[392] BLB[393] BLB[394] BLB[395]
+ GBL[98] GBLB[98] GW[98] GWB[98] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_99 BL[396] BL[397] BL[398] BL[399] BLB[396] BLB[397] BLB[398] BLB[399]
+ GBL[99] GBLB[99] GW[99] GWB[99] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_100 BL[400] BL[401] BL[402] BL[403] BLB[400] BLB[401] BLB[402] BLB[403]
+ GBL[100] GBLB[100] GW[100] GWB[100] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_101 BL[404] BL[405] BL[406] BL[407] BLB[404] BLB[405] BLB[406] BLB[407]
+ GBL[101] GBLB[101] GW[101] GWB[101] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_102 BL[408] BL[409] BL[410] BL[411] BLB[408] BLB[409] BLB[410] BLB[411]
+ GBL[102] GBLB[102] GW[102] GWB[102] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_103 BL[412] BL[413] BL[414] BL[415] BLB[412] BLB[413] BLB[414] BLB[415]
+ GBL[103] GBLB[103] GW[103] GWB[103] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_104 BL[416] BL[417] BL[418] BL[419] BLB[416] BLB[417] BLB[418] BLB[419]
+ GBL[104] GBLB[104] GW[104] GWB[104] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_105 BL[420] BL[421] BL[422] BL[423] BLB[420] BLB[421] BLB[422] BLB[423]
+ GBL[105] GBLB[105] GW[105] GWB[105] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_106 BL[424] BL[425] BL[426] BL[427] BLB[424] BLB[425] BLB[426] BLB[427]
+ GBL[106] GBLB[106] GW[106] GWB[106] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_107 BL[428] BL[429] BL[430] BL[431] BLB[428] BLB[429] BLB[430] BLB[431]
+ GBL[107] GBLB[107] GW[107] GWB[107] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_108 BL[432] BL[433] BL[434] BL[435] BLB[432] BLB[433] BLB[434] BLB[435]
+ GBL[108] GBLB[108] GW[108] GWB[108] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_109 BL[436] BL[437] BL[438] BL[439] BLB[436] BLB[437] BLB[438] BLB[439]
+ GBL[109] GBLB[109] GW[109] GWB[109] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_110 BL[440] BL[441] BL[442] BL[443] BLB[440] BLB[441] BLB[442] BLB[443]
+ GBL[110] GBLB[110] GW[110] GWB[110] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_111 BL[444] BL[445] BL[446] BL[447] BLB[444] BLB[445] BLB[446] BLB[447]
+ GBL[111] GBLB[111] GW[111] GWB[111] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_112 BL[448] BL[449] BL[450] BL[451] BLB[448] BLB[449] BLB[450] BLB[451]
+ GBL[112] GBLB[112] GW[112] GWB[112] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_113 BL[452] BL[453] BL[454] BL[455] BLB[452] BLB[453] BLB[454] BLB[455]
+ GBL[113] GBLB[113] GW[113] GWB[113] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_114 BL[456] BL[457] BL[458] BL[459] BLB[456] BLB[457] BLB[458] BLB[459]
+ GBL[114] GBLB[114] GW[114] GWB[114] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_115 BL[460] BL[461] BL[462] BL[463] BLB[460] BLB[461] BLB[462] BLB[463]
+ GBL[115] GBLB[115] GW[115] GWB[115] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_116 BL[464] BL[465] BL[466] BL[467] BLB[464] BLB[465] BLB[466] BLB[467]
+ GBL[116] GBLB[116] GW[116] GWB[116] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_117 BL[468] BL[469] BL[470] BL[471] BLB[468] BLB[469] BLB[470] BLB[471]
+ GBL[117] GBLB[117] GW[117] GWB[117] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_118 BL[472] BL[473] BL[474] BL[475] BLB[472] BLB[473] BLB[474] BLB[475]
+ GBL[118] GBLB[118] GW[118] GWB[118] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_119 BL[476] BL[477] BL[478] BL[479] BLB[476] BLB[477] BLB[478] BLB[479]
+ GBL[119] GBLB[119] GW[119] GWB[119] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_120 BL[480] BL[481] BL[482] BL[483] BLB[480] BLB[481] BLB[482] BLB[483]
+ GBL[120] GBLB[120] GW[120] GWB[120] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_121 BL[484] BL[485] BL[486] BL[487] BLB[484] BLB[485] BLB[486] BLB[487]
+ GBL[121] GBLB[121] GW[121] GWB[121] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_122 BL[488] BL[489] BL[490] BL[491] BLB[488] BLB[489] BLB[490] BLB[491]
+ GBL[122] GBLB[122] GW[122] GWB[122] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_123 BL[492] BL[493] BL[494] BL[495] BLB[492] BLB[493] BLB[494] BLB[495]
+ GBL[123] GBLB[123] GW[123] GWB[123] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_124 BL[496] BL[497] BL[498] BL[499] BLB[496] BLB[497] BLB[498] BLB[499]
+ GBL[124] GBLB[124] GW[124] GWB[124] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_125 BL[500] BL[501] BL[502] BL[503] BLB[500] BLB[501] BLB[502] BLB[503]
+ GBL[125] GBLB[125] GW[125] GWB[125] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_126 BL[504] BL[505] BL[506] BL[507] BLB[504] BLB[505] BLB[506] BLB[507]
+ GBL[126] GBLB[126] GW[126] GWB[126] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
XMCB_127 BL[508] BL[509] BL[510] BL[511] BLB[508] BLB[509] BLB[510] BLB[511]
+ GBL[127] GBLB[127] GW[127] GWB[127] VDDI VSSI WL[0] WL[1] SDBM200W80_MCB_2X4
.ENDS

.SUBCKT SDBM200W80_CELL_ARR_XY_F BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7]
+ BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18]
+ BL[19] BL[20] BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29]
+ BL[30] BL[31] BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40]
+ BL[41] BL[42] BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51]
+ BL[52] BL[53] BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62]
+ BL[63] BL[64] BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73]
+ BL[74] BL[75] BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84]
+ BL[85] BL[86] BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95]
+ BL[96] BL[97] BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105]
+ BL[106] BL[107] BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114]
+ BL[115] BL[116] BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123]
+ BL[124] BL[125] BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132]
+ BL[133] BL[134] BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141]
+ BL[142] BL[143] BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150]
+ BL[151] BL[152] BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159]
+ BL[160] BL[161] BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168]
+ BL[169] BL[170] BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177]
+ BL[178] BL[179] BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186]
+ BL[187] BL[188] BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195]
+ BL[196] BL[197] BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204]
+ BL[205] BL[206] BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213]
+ BL[214] BL[215] BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222]
+ BL[223] BL[224] BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231]
+ BL[232] BL[233] BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240]
+ BL[241] BL[242] BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249]
+ BL[250] BL[251] BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258]
+ BL[259] BL[260] BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267]
+ BL[268] BL[269] BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276]
+ BL[277] BL[278] BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285]
+ BL[286] BL[287] BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294]
+ BL[295] BL[296] BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303]
+ BL[304] BL[305] BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312]
+ BL[313] BL[314] BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321]
+ BL[322] BL[323] BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330]
+ BL[331] BL[332] BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339]
+ BL[340] BL[341] BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348]
+ BL[349] BL[350] BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357]
+ BL[358] BL[359] BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366]
+ BL[367] BL[368] BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375]
+ BL[376] BL[377] BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384]
+ BL[385] BL[386] BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393]
+ BL[394] BL[395] BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402]
+ BL[403] BL[404] BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411]
+ BL[412] BL[413] BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420]
+ BL[421] BL[422] BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429]
+ BL[430] BL[431] BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438]
+ BL[439] BL[440] BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447]
+ BL[448] BL[449] BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456]
+ BL[457] BL[458] BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465]
+ BL[466] BL[467] BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474]
+ BL[475] BL[476] BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483]
+ BL[484] BL[485] BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492]
+ BL[493] BL[494] BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501]
+ BL[502] BL[503] BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510]
+ BL[511] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9]
+ BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18]
+ BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27]
+ BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36]
+ BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45]
+ BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54]
+ BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63]
+ BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72]
+ BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81]
+ BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90]
+ BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99]
+ BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107]
+ BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115]
+ BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123]
+ BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131]
+ BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139]
+ BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147]
+ BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155]
+ BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163]
+ BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171]
+ BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179]
+ BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187]
+ BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195]
+ BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203]
+ BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211]
+ BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219]
+ BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227]
+ BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235]
+ BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243]
+ BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251]
+ BLB[252] BLB[253] BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259]
+ BLB[260] BLB[261] BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267]
+ BLB[268] BLB[269] BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275]
+ BLB[276] BLB[277] BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283]
+ BLB[284] BLB[285] BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291]
+ BLB[292] BLB[293] BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299]
+ BLB[300] BLB[301] BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307]
+ BLB[308] BLB[309] BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315]
+ BLB[316] BLB[317] BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323]
+ BLB[324] BLB[325] BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331]
+ BLB[332] BLB[333] BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339]
+ BLB[340] BLB[341] BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347]
+ BLB[348] BLB[349] BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355]
+ BLB[356] BLB[357] BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363]
+ BLB[364] BLB[365] BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371]
+ BLB[372] BLB[373] BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379]
+ BLB[380] BLB[381] BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387]
+ BLB[388] BLB[389] BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395]
+ BLB[396] BLB[397] BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403]
+ BLB[404] BLB[405] BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411]
+ BLB[412] BLB[413] BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419]
+ BLB[420] BLB[421] BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427]
+ BLB[428] BLB[429] BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435]
+ BLB[436] BLB[437] BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443]
+ BLB[444] BLB[445] BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451]
+ BLB[452] BLB[453] BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459]
+ BLB[460] BLB[461] BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467]
+ BLB[468] BLB[469] BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475]
+ BLB[476] BLB[477] BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483]
+ BLB[484] BLB[485] BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491]
+ BLB[492] BLB[493] BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499]
+ BLB[500] BLB[501] BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507]
+ BLB[508] BLB[509] BLB[510] BLB[511] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6]
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17]
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28]
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39]
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50]
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61]
+ WL[62] WL[63] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6]
+ GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16]
+ GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25]
+ GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34]
+ GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43]
+ GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52]
+ GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61]
+ GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69] GBL[70]
+ GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78] GBL[79]
+ GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87] GBL[88]
+ GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96] GBL[97]
+ GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105] GBL[106]
+ GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113] GBL[114]
+ GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121] GBL[122]
+ GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2] GBLB[3]
+ GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12]
+ GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20]
+ GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28]
+ GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36]
+ GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44]
+ GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52]
+ GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60]
+ GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67] GBLB[68]
+ GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75] GBLB[76]
+ GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83] GBLB[84]
+ GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91] GBLB[92]
+ GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99] GBLB[100]
+ GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106] GBLB[107]
+ GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113] GBLB[114]
+ GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120] GBLB[121]
+ GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0] GW[1] GW[2]
+ GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14]
+ GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25]
+ GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36]
+ GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47]
+ GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58]
+ GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67] GW[68] GW[69]
+ GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78] GW[79] GW[80]
+ GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89] GW[90] GW[91]
+ GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100] GW[101]
+ GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109] GW[110]
+ GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118] GW[119]
+ GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127]
XCELL_ARR_X_0 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[0] WL[1] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_1 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[2] WL[3] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_2 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[4] WL[5] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_3 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[6] WL[7] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_4 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[8] WL[9] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_5 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[10] WL[11] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_6 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[12] WL[13] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_7 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[14] WL[15] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_8 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[16] WL[17] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_9 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261] BLB[262]
+ BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269] BLB[270]
+ BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277] BLB[278]
+ BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285] BLB[286]
+ BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293] BLB[294]
+ BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301] BLB[302]
+ BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309] BLB[310]
+ BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317] BLB[318]
+ BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325] BLB[326]
+ BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333] BLB[334]
+ BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341] BLB[342]
+ BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349] BLB[350]
+ BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357] BLB[358]
+ BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365] BLB[366]
+ BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373] BLB[374]
+ BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381] BLB[382]
+ BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389] BLB[390]
+ BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397] BLB[398]
+ BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405] BLB[406]
+ BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413] BLB[414]
+ BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421] BLB[422]
+ BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429] BLB[430]
+ BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437] BLB[438]
+ BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445] BLB[446]
+ BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453] BLB[454]
+ BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461] BLB[462]
+ BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469] BLB[470]
+ BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477] BLB[478]
+ BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485] BLB[486]
+ BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493] BLB[494]
+ BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501] BLB[502]
+ BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509] BLB[510]
+ BLB[511] WL[18] WL[19] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69]
+ GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78]
+ GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87]
+ GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96]
+ GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105]
+ GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113]
+ GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121]
+ GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2]
+ GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11]
+ GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35]
+ GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43]
+ GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51]
+ GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_10 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[20] WL[21] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_11 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[22] WL[23] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_12 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[24] WL[25] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_13 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[26] WL[27] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_14 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[28] WL[29] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_15 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[30] WL[31] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_16 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[32] WL[33] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_17 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[34] WL[35] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_18 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[36] WL[37] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_19 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[38] WL[39] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_20 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[40] WL[41] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_21 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[42] WL[43] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_22 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[44] WL[45] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_23 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[46] WL[47] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_24 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[48] WL[49] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_25 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[50] WL[51] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_26 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[52] WL[53] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_27 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[54] WL[55] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_28 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[56] WL[57] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_29 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[58] WL[59] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_30 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[60] WL[61] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
XCELL_ARR_X_31 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] WL[62] WL[63] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41]
+ GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50]
+ GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59]
+ GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68]
+ GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77]
+ GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86]
+ GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95]
+ GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104]
+ GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112]
+ GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120]
+ GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66]
+ GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74]
+ GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82]
+ GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90]
+ GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98]
+ GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67]
+ GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78]
+ GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89]
+ GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100]
+ GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109]
+ GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118]
+ GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_X
.ENDS

.SUBCKT SDBM200W80_LIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6]
+ GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16]
+ GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25]
+ GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34]
+ GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43]
+ GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52]
+ GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61]
+ GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69] GBL[70]
+ GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78] GBL[79]
+ GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87] GBL[88]
+ GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96] GBL[97]
+ GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105] GBL[106]
+ GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113] GBL[114]
+ GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121] GBL[122]
+ GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2] GBLB[3]
+ GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12]
+ GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20]
+ GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28]
+ GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36]
+ GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44]
+ GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52]
+ GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60]
+ GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67] GBLB[68]
+ GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75] GBLB[76]
+ GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83] GBLB[84]
+ GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91] GBLB[92]
+ GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99] GBLB[100]
+ GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106] GBLB[107]
+ GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113] GBLB[114]
+ GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120] GBLB[121]
+ GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] LIOPD WL[0] WL[1]
+ WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13]
+ WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24]
+ WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35]
+ WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46]
+ WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57]
+ WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68]
+ WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79]
+ WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90]
+ WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101]
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110]
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119]
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] BLEQ_DN
+ BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10]
+ GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21]
+ GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32]
+ GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43]
+ GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54]
+ GW[55] GW[56] GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65]
+ GW[66] GW[67] GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76]
+ GW[77] GW[78] GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87]
+ GW[88] GW[89] GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98]
+ GW[99] GW[100] GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108]
+ GW[109] GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117]
+ GW[118] GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126]
+ GW[127] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9]
+ GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18]
+ GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27]
+ GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36]
+ GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45]
+ GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54]
+ GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63]
+ GWB[64] GWB[65] GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72]
+ GWB[73] GWB[74] GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81]
+ GWB[82] GWB[83] GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90]
+ GWB[91] GWB[92] GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99]
+ GWB[100] GWB[101] GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107]
+ GWB[108] GWB[109] GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115]
+ GWB[116] GWB[117] GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123]
+ GWB[124] GWB[125] GWB[126] GWB[127] PREBG SAEB Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] VDDI VSSI
XCELL_ARR_DN_F BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6]
+ BL_DN[7] BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14]
+ BL_DN[15] BL_DN[16] BL_DN[17] BL_DN[18] BL_DN[19] BL_DN[20] BL_DN[21]
+ BL_DN[22] BL_DN[23] BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27] BL_DN[28]
+ BL_DN[29] BL_DN[30] BL_DN[31] BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35]
+ BL_DN[36] BL_DN[37] BL_DN[38] BL_DN[39] BL_DN[40] BL_DN[41] BL_DN[42]
+ BL_DN[43] BL_DN[44] BL_DN[45] BL_DN[46] BL_DN[47] BL_DN[48] BL_DN[49]
+ BL_DN[50] BL_DN[51] BL_DN[52] BL_DN[53] BL_DN[54] BL_DN[55] BL_DN[56]
+ BL_DN[57] BL_DN[58] BL_DN[59] BL_DN[60] BL_DN[61] BL_DN[62] BL_DN[63]
+ BL_DN[64] BL_DN[65] BL_DN[66] BL_DN[67] BL_DN[68] BL_DN[69] BL_DN[70]
+ BL_DN[71] BL_DN[72] BL_DN[73] BL_DN[74] BL_DN[75] BL_DN[76] BL_DN[77]
+ BL_DN[78] BL_DN[79] BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83] BL_DN[84]
+ BL_DN[85] BL_DN[86] BL_DN[87] BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91]
+ BL_DN[92] BL_DN[93] BL_DN[94] BL_DN[95] BL_DN[96] BL_DN[97] BL_DN[98]
+ BL_DN[99] BL_DN[100] BL_DN[101] BL_DN[102] BL_DN[103] BL_DN[104] BL_DN[105]
+ BL_DN[106] BL_DN[107] BL_DN[108] BL_DN[109] BL_DN[110] BL_DN[111] BL_DN[112]
+ BL_DN[113] BL_DN[114] BL_DN[115] BL_DN[116] BL_DN[117] BL_DN[118] BL_DN[119]
+ BL_DN[120] BL_DN[121] BL_DN[122] BL_DN[123] BL_DN[124] BL_DN[125] BL_DN[126]
+ BL_DN[127] BL_DN[128] BL_DN[129] BL_DN[130] BL_DN[131] BL_DN[132] BL_DN[133]
+ BL_DN[134] BL_DN[135] BL_DN[136] BL_DN[137] BL_DN[138] BL_DN[139] BL_DN[140]
+ BL_DN[141] BL_DN[142] BL_DN[143] BL_DN[144] BL_DN[145] BL_DN[146] BL_DN[147]
+ BL_DN[148] BL_DN[149] BL_DN[150] BL_DN[151] BL_DN[152] BL_DN[153] BL_DN[154]
+ BL_DN[155] BL_DN[156] BL_DN[157] BL_DN[158] BL_DN[159] BL_DN[160] BL_DN[161]
+ BL_DN[162] BL_DN[163] BL_DN[164] BL_DN[165] BL_DN[166] BL_DN[167] BL_DN[168]
+ BL_DN[169] BL_DN[170] BL_DN[171] BL_DN[172] BL_DN[173] BL_DN[174] BL_DN[175]
+ BL_DN[176] BL_DN[177] BL_DN[178] BL_DN[179] BL_DN[180] BL_DN[181] BL_DN[182]
+ BL_DN[183] BL_DN[184] BL_DN[185] BL_DN[186] BL_DN[187] BL_DN[188] BL_DN[189]
+ BL_DN[190] BL_DN[191] BL_DN[192] BL_DN[193] BL_DN[194] BL_DN[195] BL_DN[196]
+ BL_DN[197] BL_DN[198] BL_DN[199] BL_DN[200] BL_DN[201] BL_DN[202] BL_DN[203]
+ BL_DN[204] BL_DN[205] BL_DN[206] BL_DN[207] BL_DN[208] BL_DN[209] BL_DN[210]
+ BL_DN[211] BL_DN[212] BL_DN[213] BL_DN[214] BL_DN[215] BL_DN[216] BL_DN[217]
+ BL_DN[218] BL_DN[219] BL_DN[220] BL_DN[221] BL_DN[222] BL_DN[223] BL_DN[224]
+ BL_DN[225] BL_DN[226] BL_DN[227] BL_DN[228] BL_DN[229] BL_DN[230] BL_DN[231]
+ BL_DN[232] BL_DN[233] BL_DN[234] BL_DN[235] BL_DN[236] BL_DN[237] BL_DN[238]
+ BL_DN[239] BL_DN[240] BL_DN[241] BL_DN[242] BL_DN[243] BL_DN[244] BL_DN[245]
+ BL_DN[246] BL_DN[247] BL_DN[248] BL_DN[249] BL_DN[250] BL_DN[251] BL_DN[252]
+ BL_DN[253] BL_DN[254] BL_DN[255] BL_DN[256] BL_DN[257] BL_DN[258] BL_DN[259]
+ BL_DN[260] BL_DN[261] BL_DN[262] BL_DN[263] BL_DN[264] BL_DN[265] BL_DN[266]
+ BL_DN[267] BL_DN[268] BL_DN[269] BL_DN[270] BL_DN[271] BL_DN[272] BL_DN[273]
+ BL_DN[274] BL_DN[275] BL_DN[276] BL_DN[277] BL_DN[278] BL_DN[279] BL_DN[280]
+ BL_DN[281] BL_DN[282] BL_DN[283] BL_DN[284] BL_DN[285] BL_DN[286] BL_DN[287]
+ BL_DN[288] BL_DN[289] BL_DN[290] BL_DN[291] BL_DN[292] BL_DN[293] BL_DN[294]
+ BL_DN[295] BL_DN[296] BL_DN[297] BL_DN[298] BL_DN[299] BL_DN[300] BL_DN[301]
+ BL_DN[302] BL_DN[303] BL_DN[304] BL_DN[305] BL_DN[306] BL_DN[307] BL_DN[308]
+ BL_DN[309] BL_DN[310] BL_DN[311] BL_DN[312] BL_DN[313] BL_DN[314] BL_DN[315]
+ BL_DN[316] BL_DN[317] BL_DN[318] BL_DN[319] BL_DN[320] BL_DN[321] BL_DN[322]
+ BL_DN[323] BL_DN[324] BL_DN[325] BL_DN[326] BL_DN[327] BL_DN[328] BL_DN[329]
+ BL_DN[330] BL_DN[331] BL_DN[332] BL_DN[333] BL_DN[334] BL_DN[335] BL_DN[336]
+ BL_DN[337] BL_DN[338] BL_DN[339] BL_DN[340] BL_DN[341] BL_DN[342] BL_DN[343]
+ BL_DN[344] BL_DN[345] BL_DN[346] BL_DN[347] BL_DN[348] BL_DN[349] BL_DN[350]
+ BL_DN[351] BL_DN[352] BL_DN[353] BL_DN[354] BL_DN[355] BL_DN[356] BL_DN[357]
+ BL_DN[358] BL_DN[359] BL_DN[360] BL_DN[361] BL_DN[362] BL_DN[363] BL_DN[364]
+ BL_DN[365] BL_DN[366] BL_DN[367] BL_DN[368] BL_DN[369] BL_DN[370] BL_DN[371]
+ BL_DN[372] BL_DN[373] BL_DN[374] BL_DN[375] BL_DN[376] BL_DN[377] BL_DN[378]
+ BL_DN[379] BL_DN[380] BL_DN[381] BL_DN[382] BL_DN[383] BL_DN[384] BL_DN[385]
+ BL_DN[386] BL_DN[387] BL_DN[388] BL_DN[389] BL_DN[390] BL_DN[391] BL_DN[392]
+ BL_DN[393] BL_DN[394] BL_DN[395] BL_DN[396] BL_DN[397] BL_DN[398] BL_DN[399]
+ BL_DN[400] BL_DN[401] BL_DN[402] BL_DN[403] BL_DN[404] BL_DN[405] BL_DN[406]
+ BL_DN[407] BL_DN[408] BL_DN[409] BL_DN[410] BL_DN[411] BL_DN[412] BL_DN[413]
+ BL_DN[414] BL_DN[415] BL_DN[416] BL_DN[417] BL_DN[418] BL_DN[419] BL_DN[420]
+ BL_DN[421] BL_DN[422] BL_DN[423] BL_DN[424] BL_DN[425] BL_DN[426] BL_DN[427]
+ BL_DN[428] BL_DN[429] BL_DN[430] BL_DN[431] BL_DN[432] BL_DN[433] BL_DN[434]
+ BL_DN[435] BL_DN[436] BL_DN[437] BL_DN[438] BL_DN[439] BL_DN[440] BL_DN[441]
+ BL_DN[442] BL_DN[443] BL_DN[444] BL_DN[445] BL_DN[446] BL_DN[447] BL_DN[448]
+ BL_DN[449] BL_DN[450] BL_DN[451] BL_DN[452] BL_DN[453] BL_DN[454] BL_DN[455]
+ BL_DN[456] BL_DN[457] BL_DN[458] BL_DN[459] BL_DN[460] BL_DN[461] BL_DN[462]
+ BL_DN[463] BL_DN[464] BL_DN[465] BL_DN[466] BL_DN[467] BL_DN[468] BL_DN[469]
+ BL_DN[470] BL_DN[471] BL_DN[472] BL_DN[473] BL_DN[474] BL_DN[475] BL_DN[476]
+ BL_DN[477] BL_DN[478] BL_DN[479] BL_DN[480] BL_DN[481] BL_DN[482] BL_DN[483]
+ BL_DN[484] BL_DN[485] BL_DN[486] BL_DN[487] BL_DN[488] BL_DN[489] BL_DN[490]
+ BL_DN[491] BL_DN[492] BL_DN[493] BL_DN[494] BL_DN[495] BL_DN[496] BL_DN[497]
+ BL_DN[498] BL_DN[499] BL_DN[500] BL_DN[501] BL_DN[502] BL_DN[503] BL_DN[504]
+ BL_DN[505] BL_DN[506] BL_DN[507] BL_DN[508] BL_DN[509] BL_DN[510] BL_DN[511]
+ BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] BLB_DN[6]
+ BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] BLB_DN[13]
+ BLB_DN[14] BLB_DN[15] BLB_DN[16] BLB_DN[17] BLB_DN[18] BLB_DN[19] BLB_DN[20]
+ BLB_DN[21] BLB_DN[22] BLB_DN[23] BLB_DN[24] BLB_DN[25] BLB_DN[26] BLB_DN[27]
+ BLB_DN[28] BLB_DN[29] BLB_DN[30] BLB_DN[31] BLB_DN[32] BLB_DN[33] BLB_DN[34]
+ BLB_DN[35] BLB_DN[36] BLB_DN[37] BLB_DN[38] BLB_DN[39] BLB_DN[40] BLB_DN[41]
+ BLB_DN[42] BLB_DN[43] BLB_DN[44] BLB_DN[45] BLB_DN[46] BLB_DN[47] BLB_DN[48]
+ BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_DN[52] BLB_DN[53] BLB_DN[54] BLB_DN[55]
+ BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59] BLB_DN[60] BLB_DN[61] BLB_DN[62]
+ BLB_DN[63] BLB_DN[64] BLB_DN[65] BLB_DN[66] BLB_DN[67] BLB_DN[68] BLB_DN[69]
+ BLB_DN[70] BLB_DN[71] BLB_DN[72] BLB_DN[73] BLB_DN[74] BLB_DN[75] BLB_DN[76]
+ BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_DN[80] BLB_DN[81] BLB_DN[82] BLB_DN[83]
+ BLB_DN[84] BLB_DN[85] BLB_DN[86] BLB_DN[87] BLB_DN[88] BLB_DN[89] BLB_DN[90]
+ BLB_DN[91] BLB_DN[92] BLB_DN[93] BLB_DN[94] BLB_DN[95] BLB_DN[96] BLB_DN[97]
+ BLB_DN[98] BLB_DN[99] BLB_DN[100] BLB_DN[101] BLB_DN[102] BLB_DN[103]
+ BLB_DN[104] BLB_DN[105] BLB_DN[106] BLB_DN[107] BLB_DN[108] BLB_DN[109]
+ BLB_DN[110] BLB_DN[111] BLB_DN[112] BLB_DN[113] BLB_DN[114] BLB_DN[115]
+ BLB_DN[116] BLB_DN[117] BLB_DN[118] BLB_DN[119] BLB_DN[120] BLB_DN[121]
+ BLB_DN[122] BLB_DN[123] BLB_DN[124] BLB_DN[125] BLB_DN[126] BLB_DN[127]
+ BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131] BLB_DN[132] BLB_DN[133]
+ BLB_DN[134] BLB_DN[135] BLB_DN[136] BLB_DN[137] BLB_DN[138] BLB_DN[139]
+ BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143] BLB_DN[144] BLB_DN[145]
+ BLB_DN[146] BLB_DN[147] BLB_DN[148] BLB_DN[149] BLB_DN[150] BLB_DN[151]
+ BLB_DN[152] BLB_DN[153] BLB_DN[154] BLB_DN[155] BLB_DN[156] BLB_DN[157]
+ BLB_DN[158] BLB_DN[159] BLB_DN[160] BLB_DN[161] BLB_DN[162] BLB_DN[163]
+ BLB_DN[164] BLB_DN[165] BLB_DN[166] BLB_DN[167] BLB_DN[168] BLB_DN[169]
+ BLB_DN[170] BLB_DN[171] BLB_DN[172] BLB_DN[173] BLB_DN[174] BLB_DN[175]
+ BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179] BLB_DN[180] BLB_DN[181]
+ BLB_DN[182] BLB_DN[183] BLB_DN[184] BLB_DN[185] BLB_DN[186] BLB_DN[187]
+ BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191] BLB_DN[192] BLB_DN[193]
+ BLB_DN[194] BLB_DN[195] BLB_DN[196] BLB_DN[197] BLB_DN[198] BLB_DN[199]
+ BLB_DN[200] BLB_DN[201] BLB_DN[202] BLB_DN[203] BLB_DN[204] BLB_DN[205]
+ BLB_DN[206] BLB_DN[207] BLB_DN[208] BLB_DN[209] BLB_DN[210] BLB_DN[211]
+ BLB_DN[212] BLB_DN[213] BLB_DN[214] BLB_DN[215] BLB_DN[216] BLB_DN[217]
+ BLB_DN[218] BLB_DN[219] BLB_DN[220] BLB_DN[221] BLB_DN[222] BLB_DN[223]
+ BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227] BLB_DN[228] BLB_DN[229]
+ BLB_DN[230] BLB_DN[231] BLB_DN[232] BLB_DN[233] BLB_DN[234] BLB_DN[235]
+ BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239] BLB_DN[240] BLB_DN[241]
+ BLB_DN[242] BLB_DN[243] BLB_DN[244] BLB_DN[245] BLB_DN[246] BLB_DN[247]
+ BLB_DN[248] BLB_DN[249] BLB_DN[250] BLB_DN[251] BLB_DN[252] BLB_DN[253]
+ BLB_DN[254] BLB_DN[255] BLB_DN[256] BLB_DN[257] BLB_DN[258] BLB_DN[259]
+ BLB_DN[260] BLB_DN[261] BLB_DN[262] BLB_DN[263] BLB_DN[264] BLB_DN[265]
+ BLB_DN[266] BLB_DN[267] BLB_DN[268] BLB_DN[269] BLB_DN[270] BLB_DN[271]
+ BLB_DN[272] BLB_DN[273] BLB_DN[274] BLB_DN[275] BLB_DN[276] BLB_DN[277]
+ BLB_DN[278] BLB_DN[279] BLB_DN[280] BLB_DN[281] BLB_DN[282] BLB_DN[283]
+ BLB_DN[284] BLB_DN[285] BLB_DN[286] BLB_DN[287] BLB_DN[288] BLB_DN[289]
+ BLB_DN[290] BLB_DN[291] BLB_DN[292] BLB_DN[293] BLB_DN[294] BLB_DN[295]
+ BLB_DN[296] BLB_DN[297] BLB_DN[298] BLB_DN[299] BLB_DN[300] BLB_DN[301]
+ BLB_DN[302] BLB_DN[303] BLB_DN[304] BLB_DN[305] BLB_DN[306] BLB_DN[307]
+ BLB_DN[308] BLB_DN[309] BLB_DN[310] BLB_DN[311] BLB_DN[312] BLB_DN[313]
+ BLB_DN[314] BLB_DN[315] BLB_DN[316] BLB_DN[317] BLB_DN[318] BLB_DN[319]
+ BLB_DN[320] BLB_DN[321] BLB_DN[322] BLB_DN[323] BLB_DN[324] BLB_DN[325]
+ BLB_DN[326] BLB_DN[327] BLB_DN[328] BLB_DN[329] BLB_DN[330] BLB_DN[331]
+ BLB_DN[332] BLB_DN[333] BLB_DN[334] BLB_DN[335] BLB_DN[336] BLB_DN[337]
+ BLB_DN[338] BLB_DN[339] BLB_DN[340] BLB_DN[341] BLB_DN[342] BLB_DN[343]
+ BLB_DN[344] BLB_DN[345] BLB_DN[346] BLB_DN[347] BLB_DN[348] BLB_DN[349]
+ BLB_DN[350] BLB_DN[351] BLB_DN[352] BLB_DN[353] BLB_DN[354] BLB_DN[355]
+ BLB_DN[356] BLB_DN[357] BLB_DN[358] BLB_DN[359] BLB_DN[360] BLB_DN[361]
+ BLB_DN[362] BLB_DN[363] BLB_DN[364] BLB_DN[365] BLB_DN[366] BLB_DN[367]
+ BLB_DN[368] BLB_DN[369] BLB_DN[370] BLB_DN[371] BLB_DN[372] BLB_DN[373]
+ BLB_DN[374] BLB_DN[375] BLB_DN[376] BLB_DN[377] BLB_DN[378] BLB_DN[379]
+ BLB_DN[380] BLB_DN[381] BLB_DN[382] BLB_DN[383] BLB_DN[384] BLB_DN[385]
+ BLB_DN[386] BLB_DN[387] BLB_DN[388] BLB_DN[389] BLB_DN[390] BLB_DN[391]
+ BLB_DN[392] BLB_DN[393] BLB_DN[394] BLB_DN[395] BLB_DN[396] BLB_DN[397]
+ BLB_DN[398] BLB_DN[399] BLB_DN[400] BLB_DN[401] BLB_DN[402] BLB_DN[403]
+ BLB_DN[404] BLB_DN[405] BLB_DN[406] BLB_DN[407] BLB_DN[408] BLB_DN[409]
+ BLB_DN[410] BLB_DN[411] BLB_DN[412] BLB_DN[413] BLB_DN[414] BLB_DN[415]
+ BLB_DN[416] BLB_DN[417] BLB_DN[418] BLB_DN[419] BLB_DN[420] BLB_DN[421]
+ BLB_DN[422] BLB_DN[423] BLB_DN[424] BLB_DN[425] BLB_DN[426] BLB_DN[427]
+ BLB_DN[428] BLB_DN[429] BLB_DN[430] BLB_DN[431] BLB_DN[432] BLB_DN[433]
+ BLB_DN[434] BLB_DN[435] BLB_DN[436] BLB_DN[437] BLB_DN[438] BLB_DN[439]
+ BLB_DN[440] BLB_DN[441] BLB_DN[442] BLB_DN[443] BLB_DN[444] BLB_DN[445]
+ BLB_DN[446] BLB_DN[447] BLB_DN[448] BLB_DN[449] BLB_DN[450] BLB_DN[451]
+ BLB_DN[452] BLB_DN[453] BLB_DN[454] BLB_DN[455] BLB_DN[456] BLB_DN[457]
+ BLB_DN[458] BLB_DN[459] BLB_DN[460] BLB_DN[461] BLB_DN[462] BLB_DN[463]
+ BLB_DN[464] BLB_DN[465] BLB_DN[466] BLB_DN[467] BLB_DN[468] BLB_DN[469]
+ BLB_DN[470] BLB_DN[471] BLB_DN[472] BLB_DN[473] BLB_DN[474] BLB_DN[475]
+ BLB_DN[476] BLB_DN[477] BLB_DN[478] BLB_DN[479] BLB_DN[480] BLB_DN[481]
+ BLB_DN[482] BLB_DN[483] BLB_DN[484] BLB_DN[485] BLB_DN[486] BLB_DN[487]
+ BLB_DN[488] BLB_DN[489] BLB_DN[490] BLB_DN[491] BLB_DN[492] BLB_DN[493]
+ BLB_DN[494] BLB_DN[495] BLB_DN[496] BLB_DN[497] BLB_DN[498] BLB_DN[499]
+ BLB_DN[500] BLB_DN[501] BLB_DN[502] BLB_DN[503] BLB_DN[504] BLB_DN[505]
+ BLB_DN[506] BLB_DN[507] BLB_DN[508] BLB_DN[509] BLB_DN[510] BLB_DN[511] WL[0]
+ WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12]
+ WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23]
+ WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34]
+ WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45]
+ WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56]
+ WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] VDDI VSSI GBL[0] GBL[1]
+ GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBL[64] GBL[65]
+ GBL[66] GBL[67] GBL[68] GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74]
+ GBL[75] GBL[76] GBL[77] GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83]
+ GBL[84] GBL[85] GBL[86] GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92]
+ GBL[93] GBL[94] GBL[95] GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101]
+ GBL[102] GBL[103] GBL[104] GBL[105] GBL[106] GBL[107] GBL[108] GBL[109]
+ GBL[110] GBL[111] GBL[112] GBL[113] GBL[114] GBL[115] GBL[116] GBL[117]
+ GBL[118] GBL[119] GBL[120] GBL[121] GBL[122] GBL[123] GBL[124] GBL[125]
+ GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6]
+ GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15]
+ GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23]
+ GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31]
+ GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39]
+ GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47]
+ GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55]
+ GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63]
+ GBLB[64] GBLB[65] GBLB[66] GBLB[67] GBLB[68] GBLB[69] GBLB[70] GBLB[71]
+ GBLB[72] GBLB[73] GBLB[74] GBLB[75] GBLB[76] GBLB[77] GBLB[78] GBLB[79]
+ GBLB[80] GBLB[81] GBLB[82] GBLB[83] GBLB[84] GBLB[85] GBLB[86] GBLB[87]
+ GBLB[88] GBLB[89] GBLB[90] GBLB[91] GBLB[92] GBLB[93] GBLB[94] GBLB[95]
+ GBLB[96] GBLB[97] GBLB[98] GBLB[99] GBLB[100] GBLB[101] GBLB[102] GBLB[103]
+ GBLB[104] GBLB[105] GBLB[106] GBLB[107] GBLB[108] GBLB[109] GBLB[110]
+ GBLB[111] GBLB[112] GBLB[113] GBLB[114] GBLB[115] GBLB[116] GBLB[117]
+ GBLB[118] GBLB[119] GBLB[120] GBLB[121] GBLB[122] GBLB[123] GBLB[124]
+ GBLB[125] GBLB[126] GBLB[127] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7]
+ GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18]
+ GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29]
+ GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39] GW[40]
+ GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50] GW[51]
+ GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60] GW[61] GW[62]
+ GW[63] GW[64] GW[65] GW[66] GW[67] GW[68] GW[69] GW[70] GW[71] GW[72] GW[73]
+ GW[74] GW[75] GW[76] GW[77] GW[78] GW[79] GW[80] GW[81] GW[82] GW[83] GW[84]
+ GW[85] GW[86] GW[87] GW[88] GW[89] GW[90] GW[91] GW[92] GW[93] GW[94] GW[95]
+ GW[96] GW[97] GW[98] GW[99] GW[100] GW[101] GW[102] GW[103] GW[104] GW[105]
+ GW[106] GW[107] GW[108] GW[109] GW[110] GW[111] GW[112] GW[113] GW[114]
+ GW[115] GW[116] GW[117] GW[118] GW[119] GW[120] GW[121] GW[122] GW[123]
+ GW[124] GW[125] GW[126] GW[127] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5]
+ GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15]
+ GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24]
+ GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33]
+ GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42]
+ GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51]
+ GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60]
+ GWB[61] GWB[62] GWB[63] GWB[64] GWB[65] GWB[66] GWB[67] GWB[68] GWB[69]
+ GWB[70] GWB[71] GWB[72] GWB[73] GWB[74] GWB[75] GWB[76] GWB[77] GWB[78]
+ GWB[79] GWB[80] GWB[81] GWB[82] GWB[83] GWB[84] GWB[85] GWB[86] GWB[87]
+ GWB[88] GWB[89] GWB[90] GWB[91] GWB[92] GWB[93] GWB[94] GWB[95] GWB[96]
+ GWB[97] GWB[98] GWB[99] GWB[100] GWB[101] GWB[102] GWB[103] GWB[104] GWB[105]
+ GWB[106] GWB[107] GWB[108] GWB[109] GWB[110] GWB[111] GWB[112] GWB[113]
+ GWB[114] GWB[115] GWB[116] GWB[117] GWB[118] GWB[119] GWB[120] GWB[121]
+ GWB[122] GWB[123] GWB[124] GWB[125] GWB[126] GWB[127] SDBM200W80_CELL_ARR_XY_F
XCELL_ARR_UP_F BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6]
+ BL_UP[7] BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14]
+ BL_UP[15] BL_UP[16] BL_UP[17] BL_UP[18] BL_UP[19] BL_UP[20] BL_UP[21]
+ BL_UP[22] BL_UP[23] BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27] BL_UP[28]
+ BL_UP[29] BL_UP[30] BL_UP[31] BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35]
+ BL_UP[36] BL_UP[37] BL_UP[38] BL_UP[39] BL_UP[40] BL_UP[41] BL_UP[42]
+ BL_UP[43] BL_UP[44] BL_UP[45] BL_UP[46] BL_UP[47] BL_UP[48] BL_UP[49]
+ BL_UP[50] BL_UP[51] BL_UP[52] BL_UP[53] BL_UP[54] BL_UP[55] BL_UP[56]
+ BL_UP[57] BL_UP[58] BL_UP[59] BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63]
+ BL_UP[64] BL_UP[65] BL_UP[66] BL_UP[67] BL_UP[68] BL_UP[69] BL_UP[70]
+ BL_UP[71] BL_UP[72] BL_UP[73] BL_UP[74] BL_UP[75] BL_UP[76] BL_UP[77]
+ BL_UP[78] BL_UP[79] BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] BL_UP[84]
+ BL_UP[85] BL_UP[86] BL_UP[87] BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91]
+ BL_UP[92] BL_UP[93] BL_UP[94] BL_UP[95] BL_UP[96] BL_UP[97] BL_UP[98]
+ BL_UP[99] BL_UP[100] BL_UP[101] BL_UP[102] BL_UP[103] BL_UP[104] BL_UP[105]
+ BL_UP[106] BL_UP[107] BL_UP[108] BL_UP[109] BL_UP[110] BL_UP[111] BL_UP[112]
+ BL_UP[113] BL_UP[114] BL_UP[115] BL_UP[116] BL_UP[117] BL_UP[118] BL_UP[119]
+ BL_UP[120] BL_UP[121] BL_UP[122] BL_UP[123] BL_UP[124] BL_UP[125] BL_UP[126]
+ BL_UP[127] BL_UP[128] BL_UP[129] BL_UP[130] BL_UP[131] BL_UP[132] BL_UP[133]
+ BL_UP[134] BL_UP[135] BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] BL_UP[140]
+ BL_UP[141] BL_UP[142] BL_UP[143] BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147]
+ BL_UP[148] BL_UP[149] BL_UP[150] BL_UP[151] BL_UP[152] BL_UP[153] BL_UP[154]
+ BL_UP[155] BL_UP[156] BL_UP[157] BL_UP[158] BL_UP[159] BL_UP[160] BL_UP[161]
+ BL_UP[162] BL_UP[163] BL_UP[164] BL_UP[165] BL_UP[166] BL_UP[167] BL_UP[168]
+ BL_UP[169] BL_UP[170] BL_UP[171] BL_UP[172] BL_UP[173] BL_UP[174] BL_UP[175]
+ BL_UP[176] BL_UP[177] BL_UP[178] BL_UP[179] BL_UP[180] BL_UP[181] BL_UP[182]
+ BL_UP[183] BL_UP[184] BL_UP[185] BL_UP[186] BL_UP[187] BL_UP[188] BL_UP[189]
+ BL_UP[190] BL_UP[191] BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] BL_UP[196]
+ BL_UP[197] BL_UP[198] BL_UP[199] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203]
+ BL_UP[204] BL_UP[205] BL_UP[206] BL_UP[207] BL_UP[208] BL_UP[209] BL_UP[210]
+ BL_UP[211] BL_UP[212] BL_UP[213] BL_UP[214] BL_UP[215] BL_UP[216] BL_UP[217]
+ BL_UP[218] BL_UP[219] BL_UP[220] BL_UP[221] BL_UP[222] BL_UP[223] BL_UP[224]
+ BL_UP[225] BL_UP[226] BL_UP[227] BL_UP[228] BL_UP[229] BL_UP[230] BL_UP[231]
+ BL_UP[232] BL_UP[233] BL_UP[234] BL_UP[235] BL_UP[236] BL_UP[237] BL_UP[238]
+ BL_UP[239] BL_UP[240] BL_UP[241] BL_UP[242] BL_UP[243] BL_UP[244] BL_UP[245]
+ BL_UP[246] BL_UP[247] BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] BL_UP[252]
+ BL_UP[253] BL_UP[254] BL_UP[255] BL_UP[256] BL_UP[257] BL_UP[258] BL_UP[259]
+ BL_UP[260] BL_UP[261] BL_UP[262] BL_UP[263] BL_UP[264] BL_UP[265] BL_UP[266]
+ BL_UP[267] BL_UP[268] BL_UP[269] BL_UP[270] BL_UP[271] BL_UP[272] BL_UP[273]
+ BL_UP[274] BL_UP[275] BL_UP[276] BL_UP[277] BL_UP[278] BL_UP[279] BL_UP[280]
+ BL_UP[281] BL_UP[282] BL_UP[283] BL_UP[284] BL_UP[285] BL_UP[286] BL_UP[287]
+ BL_UP[288] BL_UP[289] BL_UP[290] BL_UP[291] BL_UP[292] BL_UP[293] BL_UP[294]
+ BL_UP[295] BL_UP[296] BL_UP[297] BL_UP[298] BL_UP[299] BL_UP[300] BL_UP[301]
+ BL_UP[302] BL_UP[303] BL_UP[304] BL_UP[305] BL_UP[306] BL_UP[307] BL_UP[308]
+ BL_UP[309] BL_UP[310] BL_UP[311] BL_UP[312] BL_UP[313] BL_UP[314] BL_UP[315]
+ BL_UP[316] BL_UP[317] BL_UP[318] BL_UP[319] BL_UP[320] BL_UP[321] BL_UP[322]
+ BL_UP[323] BL_UP[324] BL_UP[325] BL_UP[326] BL_UP[327] BL_UP[328] BL_UP[329]
+ BL_UP[330] BL_UP[331] BL_UP[332] BL_UP[333] BL_UP[334] BL_UP[335] BL_UP[336]
+ BL_UP[337] BL_UP[338] BL_UP[339] BL_UP[340] BL_UP[341] BL_UP[342] BL_UP[343]
+ BL_UP[344] BL_UP[345] BL_UP[346] BL_UP[347] BL_UP[348] BL_UP[349] BL_UP[350]
+ BL_UP[351] BL_UP[352] BL_UP[353] BL_UP[354] BL_UP[355] BL_UP[356] BL_UP[357]
+ BL_UP[358] BL_UP[359] BL_UP[360] BL_UP[361] BL_UP[362] BL_UP[363] BL_UP[364]
+ BL_UP[365] BL_UP[366] BL_UP[367] BL_UP[368] BL_UP[369] BL_UP[370] BL_UP[371]
+ BL_UP[372] BL_UP[373] BL_UP[374] BL_UP[375] BL_UP[376] BL_UP[377] BL_UP[378]
+ BL_UP[379] BL_UP[380] BL_UP[381] BL_UP[382] BL_UP[383] BL_UP[384] BL_UP[385]
+ BL_UP[386] BL_UP[387] BL_UP[388] BL_UP[389] BL_UP[390] BL_UP[391] BL_UP[392]
+ BL_UP[393] BL_UP[394] BL_UP[395] BL_UP[396] BL_UP[397] BL_UP[398] BL_UP[399]
+ BL_UP[400] BL_UP[401] BL_UP[402] BL_UP[403] BL_UP[404] BL_UP[405] BL_UP[406]
+ BL_UP[407] BL_UP[408] BL_UP[409] BL_UP[410] BL_UP[411] BL_UP[412] BL_UP[413]
+ BL_UP[414] BL_UP[415] BL_UP[416] BL_UP[417] BL_UP[418] BL_UP[419] BL_UP[420]
+ BL_UP[421] BL_UP[422] BL_UP[423] BL_UP[424] BL_UP[425] BL_UP[426] BL_UP[427]
+ BL_UP[428] BL_UP[429] BL_UP[430] BL_UP[431] BL_UP[432] BL_UP[433] BL_UP[434]
+ BL_UP[435] BL_UP[436] BL_UP[437] BL_UP[438] BL_UP[439] BL_UP[440] BL_UP[441]
+ BL_UP[442] BL_UP[443] BL_UP[444] BL_UP[445] BL_UP[446] BL_UP[447] BL_UP[448]
+ BL_UP[449] BL_UP[450] BL_UP[451] BL_UP[452] BL_UP[453] BL_UP[454] BL_UP[455]
+ BL_UP[456] BL_UP[457] BL_UP[458] BL_UP[459] BL_UP[460] BL_UP[461] BL_UP[462]
+ BL_UP[463] BL_UP[464] BL_UP[465] BL_UP[466] BL_UP[467] BL_UP[468] BL_UP[469]
+ BL_UP[470] BL_UP[471] BL_UP[472] BL_UP[473] BL_UP[474] BL_UP[475] BL_UP[476]
+ BL_UP[477] BL_UP[478] BL_UP[479] BL_UP[480] BL_UP[481] BL_UP[482] BL_UP[483]
+ BL_UP[484] BL_UP[485] BL_UP[486] BL_UP[487] BL_UP[488] BL_UP[489] BL_UP[490]
+ BL_UP[491] BL_UP[492] BL_UP[493] BL_UP[494] BL_UP[495] BL_UP[496] BL_UP[497]
+ BL_UP[498] BL_UP[499] BL_UP[500] BL_UP[501] BL_UP[502] BL_UP[503] BL_UP[504]
+ BL_UP[505] BL_UP[506] BL_UP[507] BL_UP[508] BL_UP[509] BL_UP[510] BL_UP[511]
+ BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] BLB_UP[5] BLB_UP[6]
+ BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] BLB_UP[11] BLB_UP[12] BLB_UP[13]
+ BLB_UP[14] BLB_UP[15] BLB_UP[16] BLB_UP[17] BLB_UP[18] BLB_UP[19] BLB_UP[20]
+ BLB_UP[21] BLB_UP[22] BLB_UP[23] BLB_UP[24] BLB_UP[25] BLB_UP[26] BLB_UP[27]
+ BLB_UP[28] BLB_UP[29] BLB_UP[30] BLB_UP[31] BLB_UP[32] BLB_UP[33] BLB_UP[34]
+ BLB_UP[35] BLB_UP[36] BLB_UP[37] BLB_UP[38] BLB_UP[39] BLB_UP[40] BLB_UP[41]
+ BLB_UP[42] BLB_UP[43] BLB_UP[44] BLB_UP[45] BLB_UP[46] BLB_UP[47] BLB_UP[48]
+ BLB_UP[49] BLB_UP[50] BLB_UP[51] BLB_UP[52] BLB_UP[53] BLB_UP[54] BLB_UP[55]
+ BLB_UP[56] BLB_UP[57] BLB_UP[58] BLB_UP[59] BLB_UP[60] BLB_UP[61] BLB_UP[62]
+ BLB_UP[63] BLB_UP[64] BLB_UP[65] BLB_UP[66] BLB_UP[67] BLB_UP[68] BLB_UP[69]
+ BLB_UP[70] BLB_UP[71] BLB_UP[72] BLB_UP[73] BLB_UP[74] BLB_UP[75] BLB_UP[76]
+ BLB_UP[77] BLB_UP[78] BLB_UP[79] BLB_UP[80] BLB_UP[81] BLB_UP[82] BLB_UP[83]
+ BLB_UP[84] BLB_UP[85] BLB_UP[86] BLB_UP[87] BLB_UP[88] BLB_UP[89] BLB_UP[90]
+ BLB_UP[91] BLB_UP[92] BLB_UP[93] BLB_UP[94] BLB_UP[95] BLB_UP[96] BLB_UP[97]
+ BLB_UP[98] BLB_UP[99] BLB_UP[100] BLB_UP[101] BLB_UP[102] BLB_UP[103]
+ BLB_UP[104] BLB_UP[105] BLB_UP[106] BLB_UP[107] BLB_UP[108] BLB_UP[109]
+ BLB_UP[110] BLB_UP[111] BLB_UP[112] BLB_UP[113] BLB_UP[114] BLB_UP[115]
+ BLB_UP[116] BLB_UP[117] BLB_UP[118] BLB_UP[119] BLB_UP[120] BLB_UP[121]
+ BLB_UP[122] BLB_UP[123] BLB_UP[124] BLB_UP[125] BLB_UP[126] BLB_UP[127]
+ BLB_UP[128] BLB_UP[129] BLB_UP[130] BLB_UP[131] BLB_UP[132] BLB_UP[133]
+ BLB_UP[134] BLB_UP[135] BLB_UP[136] BLB_UP[137] BLB_UP[138] BLB_UP[139]
+ BLB_UP[140] BLB_UP[141] BLB_UP[142] BLB_UP[143] BLB_UP[144] BLB_UP[145]
+ BLB_UP[146] BLB_UP[147] BLB_UP[148] BLB_UP[149] BLB_UP[150] BLB_UP[151]
+ BLB_UP[152] BLB_UP[153] BLB_UP[154] BLB_UP[155] BLB_UP[156] BLB_UP[157]
+ BLB_UP[158] BLB_UP[159] BLB_UP[160] BLB_UP[161] BLB_UP[162] BLB_UP[163]
+ BLB_UP[164] BLB_UP[165] BLB_UP[166] BLB_UP[167] BLB_UP[168] BLB_UP[169]
+ BLB_UP[170] BLB_UP[171] BLB_UP[172] BLB_UP[173] BLB_UP[174] BLB_UP[175]
+ BLB_UP[176] BLB_UP[177] BLB_UP[178] BLB_UP[179] BLB_UP[180] BLB_UP[181]
+ BLB_UP[182] BLB_UP[183] BLB_UP[184] BLB_UP[185] BLB_UP[186] BLB_UP[187]
+ BLB_UP[188] BLB_UP[189] BLB_UP[190] BLB_UP[191] BLB_UP[192] BLB_UP[193]
+ BLB_UP[194] BLB_UP[195] BLB_UP[196] BLB_UP[197] BLB_UP[198] BLB_UP[199]
+ BLB_UP[200] BLB_UP[201] BLB_UP[202] BLB_UP[203] BLB_UP[204] BLB_UP[205]
+ BLB_UP[206] BLB_UP[207] BLB_UP[208] BLB_UP[209] BLB_UP[210] BLB_UP[211]
+ BLB_UP[212] BLB_UP[213] BLB_UP[214] BLB_UP[215] BLB_UP[216] BLB_UP[217]
+ BLB_UP[218] BLB_UP[219] BLB_UP[220] BLB_UP[221] BLB_UP[222] BLB_UP[223]
+ BLB_UP[224] BLB_UP[225] BLB_UP[226] BLB_UP[227] BLB_UP[228] BLB_UP[229]
+ BLB_UP[230] BLB_UP[231] BLB_UP[232] BLB_UP[233] BLB_UP[234] BLB_UP[235]
+ BLB_UP[236] BLB_UP[237] BLB_UP[238] BLB_UP[239] BLB_UP[240] BLB_UP[241]
+ BLB_UP[242] BLB_UP[243] BLB_UP[244] BLB_UP[245] BLB_UP[246] BLB_UP[247]
+ BLB_UP[248] BLB_UP[249] BLB_UP[250] BLB_UP[251] BLB_UP[252] BLB_UP[253]
+ BLB_UP[254] BLB_UP[255] BLB_UP[256] BLB_UP[257] BLB_UP[258] BLB_UP[259]
+ BLB_UP[260] BLB_UP[261] BLB_UP[262] BLB_UP[263] BLB_UP[264] BLB_UP[265]
+ BLB_UP[266] BLB_UP[267] BLB_UP[268] BLB_UP[269] BLB_UP[270] BLB_UP[271]
+ BLB_UP[272] BLB_UP[273] BLB_UP[274] BLB_UP[275] BLB_UP[276] BLB_UP[277]
+ BLB_UP[278] BLB_UP[279] BLB_UP[280] BLB_UP[281] BLB_UP[282] BLB_UP[283]
+ BLB_UP[284] BLB_UP[285] BLB_UP[286] BLB_UP[287] BLB_UP[288] BLB_UP[289]
+ BLB_UP[290] BLB_UP[291] BLB_UP[292] BLB_UP[293] BLB_UP[294] BLB_UP[295]
+ BLB_UP[296] BLB_UP[297] BLB_UP[298] BLB_UP[299] BLB_UP[300] BLB_UP[301]
+ BLB_UP[302] BLB_UP[303] BLB_UP[304] BLB_UP[305] BLB_UP[306] BLB_UP[307]
+ BLB_UP[308] BLB_UP[309] BLB_UP[310] BLB_UP[311] BLB_UP[312] BLB_UP[313]
+ BLB_UP[314] BLB_UP[315] BLB_UP[316] BLB_UP[317] BLB_UP[318] BLB_UP[319]
+ BLB_UP[320] BLB_UP[321] BLB_UP[322] BLB_UP[323] BLB_UP[324] BLB_UP[325]
+ BLB_UP[326] BLB_UP[327] BLB_UP[328] BLB_UP[329] BLB_UP[330] BLB_UP[331]
+ BLB_UP[332] BLB_UP[333] BLB_UP[334] BLB_UP[335] BLB_UP[336] BLB_UP[337]
+ BLB_UP[338] BLB_UP[339] BLB_UP[340] BLB_UP[341] BLB_UP[342] BLB_UP[343]
+ BLB_UP[344] BLB_UP[345] BLB_UP[346] BLB_UP[347] BLB_UP[348] BLB_UP[349]
+ BLB_UP[350] BLB_UP[351] BLB_UP[352] BLB_UP[353] BLB_UP[354] BLB_UP[355]
+ BLB_UP[356] BLB_UP[357] BLB_UP[358] BLB_UP[359] BLB_UP[360] BLB_UP[361]
+ BLB_UP[362] BLB_UP[363] BLB_UP[364] BLB_UP[365] BLB_UP[366] BLB_UP[367]
+ BLB_UP[368] BLB_UP[369] BLB_UP[370] BLB_UP[371] BLB_UP[372] BLB_UP[373]
+ BLB_UP[374] BLB_UP[375] BLB_UP[376] BLB_UP[377] BLB_UP[378] BLB_UP[379]
+ BLB_UP[380] BLB_UP[381] BLB_UP[382] BLB_UP[383] BLB_UP[384] BLB_UP[385]
+ BLB_UP[386] BLB_UP[387] BLB_UP[388] BLB_UP[389] BLB_UP[390] BLB_UP[391]
+ BLB_UP[392] BLB_UP[393] BLB_UP[394] BLB_UP[395] BLB_UP[396] BLB_UP[397]
+ BLB_UP[398] BLB_UP[399] BLB_UP[400] BLB_UP[401] BLB_UP[402] BLB_UP[403]
+ BLB_UP[404] BLB_UP[405] BLB_UP[406] BLB_UP[407] BLB_UP[408] BLB_UP[409]
+ BLB_UP[410] BLB_UP[411] BLB_UP[412] BLB_UP[413] BLB_UP[414] BLB_UP[415]
+ BLB_UP[416] BLB_UP[417] BLB_UP[418] BLB_UP[419] BLB_UP[420] BLB_UP[421]
+ BLB_UP[422] BLB_UP[423] BLB_UP[424] BLB_UP[425] BLB_UP[426] BLB_UP[427]
+ BLB_UP[428] BLB_UP[429] BLB_UP[430] BLB_UP[431] BLB_UP[432] BLB_UP[433]
+ BLB_UP[434] BLB_UP[435] BLB_UP[436] BLB_UP[437] BLB_UP[438] BLB_UP[439]
+ BLB_UP[440] BLB_UP[441] BLB_UP[442] BLB_UP[443] BLB_UP[444] BLB_UP[445]
+ BLB_UP[446] BLB_UP[447] BLB_UP[448] BLB_UP[449] BLB_UP[450] BLB_UP[451]
+ BLB_UP[452] BLB_UP[453] BLB_UP[454] BLB_UP[455] BLB_UP[456] BLB_UP[457]
+ BLB_UP[458] BLB_UP[459] BLB_UP[460] BLB_UP[461] BLB_UP[462] BLB_UP[463]
+ BLB_UP[464] BLB_UP[465] BLB_UP[466] BLB_UP[467] BLB_UP[468] BLB_UP[469]
+ BLB_UP[470] BLB_UP[471] BLB_UP[472] BLB_UP[473] BLB_UP[474] BLB_UP[475]
+ BLB_UP[476] BLB_UP[477] BLB_UP[478] BLB_UP[479] BLB_UP[480] BLB_UP[481]
+ BLB_UP[482] BLB_UP[483] BLB_UP[484] BLB_UP[485] BLB_UP[486] BLB_UP[487]
+ BLB_UP[488] BLB_UP[489] BLB_UP[490] BLB_UP[491] BLB_UP[492] BLB_UP[493]
+ BLB_UP[494] BLB_UP[495] BLB_UP[496] BLB_UP[497] BLB_UP[498] BLB_UP[499]
+ BLB_UP[500] BLB_UP[501] BLB_UP[502] BLB_UP[503] BLB_UP[504] BLB_UP[505]
+ BLB_UP[506] BLB_UP[507] BLB_UP[508] BLB_UP[509] BLB_UP[510] BLB_UP[511] WL[64]
+ WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75]
+ WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86]
+ WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97]
+ WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107]
+ WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116]
+ WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125]
+ WL[126] WL[127] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6]
+ GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16]
+ GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25]
+ GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34]
+ GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43]
+ GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52]
+ GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61]
+ GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69] GBL[70]
+ GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78] GBL[79]
+ GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87] GBL[88]
+ GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96] GBL[97]
+ GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105] GBL[106]
+ GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113] GBL[114]
+ GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121] GBL[122]
+ GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2] GBLB[3]
+ GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12]
+ GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20]
+ GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28]
+ GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36]
+ GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44]
+ GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52]
+ GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60]
+ GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67] GBLB[68]
+ GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75] GBLB[76]
+ GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83] GBLB[84]
+ GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91] GBLB[92]
+ GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99] GBLB[100]
+ GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106] GBLB[107]
+ GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113] GBLB[114]
+ GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120] GBLB[121]
+ GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0] GW[1] GW[2]
+ GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14]
+ GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25]
+ GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36]
+ GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47]
+ GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58]
+ GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67] GW[68] GW[69]
+ GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78] GW[79] GW[80]
+ GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89] GW[90] GW[91]
+ GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100] GW[101]
+ GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109] GW[110]
+ GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118] GW[119]
+ GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SDBM200W80_CELL_ARR_XY_F
XLIO_M4_0 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_UP[0] BLB_UP[1] BLB_UP[2]
+ BLB_UP[3] BLEQ_DN BLEQ_UP BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_UP[0]
+ BL_UP[1] BL_UP[2] BL_UP[3] GBL[0] GBLB[0] GW[0] GWB[0] PREBG SAEB VDDI VSSI
+ Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0]
+ Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_1 BLB_DN[4] BLB_DN[5] BLB_DN[6] BLB_DN[7] BLB_UP[4] BLB_UP[5] BLB_UP[6]
+ BLB_UP[7] BLEQ_DN BLEQ_UP BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] BL_UP[4]
+ BL_UP[5] BL_UP[6] BL_UP[7] GBL[1] GBLB[1] GW[1] GWB[1] PREBG SAEB VDDI VSSI
+ Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0]
+ Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_2 BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_UP[8] BLB_UP[9]
+ BLB_UP[10] BLB_UP[11] BLEQ_DN BLEQ_UP BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11]
+ BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] GBL[2] GBLB[2] GW[2] GWB[2] PREBG SAEB
+ VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_3 BLB_DN[12] BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_UP[12] BLB_UP[13]
+ BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP BL_DN[12] BL_DN[13] BL_DN[14] BL_DN[15]
+ BL_UP[12] BL_UP[13] BL_UP[14] BL_UP[15] GBL[3] GBLB[3] GW[3] GWB[3] PREBG SAEB
+ VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_4 BLB_DN[16] BLB_DN[17] BLB_DN[18] BLB_DN[19] BLB_UP[16] BLB_UP[17]
+ BLB_UP[18] BLB_UP[19] BLEQ_DN BLEQ_UP BL_DN[16] BL_DN[17] BL_DN[18] BL_DN[19]
+ BL_UP[16] BL_UP[17] BL_UP[18] BL_UP[19] GBL[4] GBLB[4] GW[4] GWB[4] PREBG SAEB
+ VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_5 BLB_DN[20] BLB_DN[21] BLB_DN[22] BLB_DN[23] BLB_UP[20] BLB_UP[21]
+ BLB_UP[22] BLB_UP[23] BLEQ_DN BLEQ_UP BL_DN[20] BL_DN[21] BL_DN[22] BL_DN[23]
+ BL_UP[20] BL_UP[21] BL_UP[22] BL_UP[23] GBL[5] GBLB[5] GW[5] GWB[5] PREBG SAEB
+ VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_6 BLB_DN[24] BLB_DN[25] BLB_DN[26] BLB_DN[27] BLB_UP[24] BLB_UP[25]
+ BLB_UP[26] BLB_UP[27] BLEQ_DN BLEQ_UP BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27]
+ BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27] GBL[6] GBLB[6] GW[6] GWB[6] PREBG SAEB
+ VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_7 BLB_DN[28] BLB_DN[29] BLB_DN[30] BLB_DN[31] BLB_UP[28] BLB_UP[29]
+ BLB_UP[30] BLB_UP[31] BLEQ_DN BLEQ_UP BL_DN[28] BL_DN[29] BL_DN[30] BL_DN[31]
+ BL_UP[28] BL_UP[29] BL_UP[30] BL_UP[31] GBL[7] GBLB[7] GW[7] GWB[7] PREBG SAEB
+ VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_8 BLB_DN[32] BLB_DN[33] BLB_DN[34] BLB_DN[35] BLB_UP[32] BLB_UP[33]
+ BLB_UP[34] BLB_UP[35] BLEQ_DN BLEQ_UP BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35]
+ BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35] GBL[8] GBLB[8] GW[8] GWB[8] PREBG SAEB
+ VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_9 BLB_DN[36] BLB_DN[37] BLB_DN[38] BLB_DN[39] BLB_UP[36] BLB_UP[37]
+ BLB_UP[38] BLB_UP[39] BLEQ_DN BLEQ_UP BL_DN[36] BL_DN[37] BL_DN[38] BL_DN[39]
+ BL_UP[36] BL_UP[37] BL_UP[38] BL_UP[39] GBL[9] GBLB[9] GW[9] GWB[9] PREBG SAEB
+ VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_10 BLB_DN[40] BLB_DN[41] BLB_DN[42] BLB_DN[43] BLB_UP[40] BLB_UP[41]
+ BLB_UP[42] BLB_UP[43] BLEQ_DN BLEQ_UP BL_DN[40] BL_DN[41] BL_DN[42] BL_DN[43]
+ BL_UP[40] BL_UP[41] BL_UP[42] BL_UP[43] GBL[10] GBLB[10] GW[10] GWB[10] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_11 BLB_DN[44] BLB_DN[45] BLB_DN[46] BLB_DN[47] BLB_UP[44] BLB_UP[45]
+ BLB_UP[46] BLB_UP[47] BLEQ_DN BLEQ_UP BL_DN[44] BL_DN[45] BL_DN[46] BL_DN[47]
+ BL_UP[44] BL_UP[45] BL_UP[46] BL_UP[47] GBL[11] GBLB[11] GW[11] GWB[11] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_12 BLB_DN[48] BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_UP[48] BLB_UP[49]
+ BLB_UP[50] BLB_UP[51] BLEQ_DN BLEQ_UP BL_DN[48] BL_DN[49] BL_DN[50] BL_DN[51]
+ BL_UP[48] BL_UP[49] BL_UP[50] BL_UP[51] GBL[12] GBLB[12] GW[12] GWB[12] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_13 BLB_DN[52] BLB_DN[53] BLB_DN[54] BLB_DN[55] BLB_UP[52] BLB_UP[53]
+ BLB_UP[54] BLB_UP[55] BLEQ_DN BLEQ_UP BL_DN[52] BL_DN[53] BL_DN[54] BL_DN[55]
+ BL_UP[52] BL_UP[53] BL_UP[54] BL_UP[55] GBL[13] GBLB[13] GW[13] GWB[13] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_14 BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59] BLB_UP[56] BLB_UP[57]
+ BLB_UP[58] BLB_UP[59] BLEQ_DN BLEQ_UP BL_DN[56] BL_DN[57] BL_DN[58] BL_DN[59]
+ BL_UP[56] BL_UP[57] BL_UP[58] BL_UP[59] GBL[14] GBLB[14] GW[14] GWB[14] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_15 BLB_DN[60] BLB_DN[61] BLB_DN[62] BLB_DN[63] BLB_UP[60] BLB_UP[61]
+ BLB_UP[62] BLB_UP[63] BLEQ_DN BLEQ_UP BL_DN[60] BL_DN[61] BL_DN[62] BL_DN[63]
+ BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63] GBL[15] GBLB[15] GW[15] GWB[15] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_16 BLB_DN[64] BLB_DN[65] BLB_DN[66] BLB_DN[67] BLB_UP[64] BLB_UP[65]
+ BLB_UP[66] BLB_UP[67] BLEQ_DN BLEQ_UP BL_DN[64] BL_DN[65] BL_DN[66] BL_DN[67]
+ BL_UP[64] BL_UP[65] BL_UP[66] BL_UP[67] GBL[16] GBLB[16] GW[16] GWB[16] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_17 BLB_DN[68] BLB_DN[69] BLB_DN[70] BLB_DN[71] BLB_UP[68] BLB_UP[69]
+ BLB_UP[70] BLB_UP[71] BLEQ_DN BLEQ_UP BL_DN[68] BL_DN[69] BL_DN[70] BL_DN[71]
+ BL_UP[68] BL_UP[69] BL_UP[70] BL_UP[71] GBL[17] GBLB[17] GW[17] GWB[17] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_18 BLB_DN[72] BLB_DN[73] BLB_DN[74] BLB_DN[75] BLB_UP[72] BLB_UP[73]
+ BLB_UP[74] BLB_UP[75] BLEQ_DN BLEQ_UP BL_DN[72] BL_DN[73] BL_DN[74] BL_DN[75]
+ BL_UP[72] BL_UP[73] BL_UP[74] BL_UP[75] GBL[18] GBLB[18] GW[18] GWB[18] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_19 BLB_DN[76] BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_UP[76] BLB_UP[77]
+ BLB_UP[78] BLB_UP[79] BLEQ_DN BLEQ_UP BL_DN[76] BL_DN[77] BL_DN[78] BL_DN[79]
+ BL_UP[76] BL_UP[77] BL_UP[78] BL_UP[79] GBL[19] GBLB[19] GW[19] GWB[19] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_20 BLB_DN[80] BLB_DN[81] BLB_DN[82] BLB_DN[83] BLB_UP[80] BLB_UP[81]
+ BLB_UP[82] BLB_UP[83] BLEQ_DN BLEQ_UP BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83]
+ BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] GBL[20] GBLB[20] GW[20] GWB[20] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_21 BLB_DN[84] BLB_DN[85] BLB_DN[86] BLB_DN[87] BLB_UP[84] BLB_UP[85]
+ BLB_UP[86] BLB_UP[87] BLEQ_DN BLEQ_UP BL_DN[84] BL_DN[85] BL_DN[86] BL_DN[87]
+ BL_UP[84] BL_UP[85] BL_UP[86] BL_UP[87] GBL[21] GBLB[21] GW[21] GWB[21] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_22 BLB_DN[88] BLB_DN[89] BLB_DN[90] BLB_DN[91] BLB_UP[88] BLB_UP[89]
+ BLB_UP[90] BLB_UP[91] BLEQ_DN BLEQ_UP BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91]
+ BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91] GBL[22] GBLB[22] GW[22] GWB[22] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_23 BLB_DN[92] BLB_DN[93] BLB_DN[94] BLB_DN[95] BLB_UP[92] BLB_UP[93]
+ BLB_UP[94] BLB_UP[95] BLEQ_DN BLEQ_UP BL_DN[92] BL_DN[93] BL_DN[94] BL_DN[95]
+ BL_UP[92] BL_UP[93] BL_UP[94] BL_UP[95] GBL[23] GBLB[23] GW[23] GWB[23] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_24 BLB_DN[96] BLB_DN[97] BLB_DN[98] BLB_DN[99] BLB_UP[96] BLB_UP[97]
+ BLB_UP[98] BLB_UP[99] BLEQ_DN BLEQ_UP BL_DN[96] BL_DN[97] BL_DN[98] BL_DN[99]
+ BL_UP[96] BL_UP[97] BL_UP[98] BL_UP[99] GBL[24] GBLB[24] GW[24] GWB[24] PREBG
+ SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ SDBM200W80_LIO_M4
XLIO_M4_25 BLB_DN[100] BLB_DN[101] BLB_DN[102] BLB_DN[103] BLB_UP[100]
+ BLB_UP[101] BLB_UP[102] BLB_UP[103] BLEQ_DN BLEQ_UP BL_DN[100] BL_DN[101]
+ BL_DN[102] BL_DN[103] BL_UP[100] BL_UP[101] BL_UP[102] BL_UP[103] GBL[25]
+ GBLB[25] GW[25] GWB[25] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_26 BLB_DN[104] BLB_DN[105] BLB_DN[106] BLB_DN[107] BLB_UP[104]
+ BLB_UP[105] BLB_UP[106] BLB_UP[107] BLEQ_DN BLEQ_UP BL_DN[104] BL_DN[105]
+ BL_DN[106] BL_DN[107] BL_UP[104] BL_UP[105] BL_UP[106] BL_UP[107] GBL[26]
+ GBLB[26] GW[26] GWB[26] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_27 BLB_DN[108] BLB_DN[109] BLB_DN[110] BLB_DN[111] BLB_UP[108]
+ BLB_UP[109] BLB_UP[110] BLB_UP[111] BLEQ_DN BLEQ_UP BL_DN[108] BL_DN[109]
+ BL_DN[110] BL_DN[111] BL_UP[108] BL_UP[109] BL_UP[110] BL_UP[111] GBL[27]
+ GBLB[27] GW[27] GWB[27] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_28 BLB_DN[112] BLB_DN[113] BLB_DN[114] BLB_DN[115] BLB_UP[112]
+ BLB_UP[113] BLB_UP[114] BLB_UP[115] BLEQ_DN BLEQ_UP BL_DN[112] BL_DN[113]
+ BL_DN[114] BL_DN[115] BL_UP[112] BL_UP[113] BL_UP[114] BL_UP[115] GBL[28]
+ GBLB[28] GW[28] GWB[28] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_29 BLB_DN[116] BLB_DN[117] BLB_DN[118] BLB_DN[119] BLB_UP[116]
+ BLB_UP[117] BLB_UP[118] BLB_UP[119] BLEQ_DN BLEQ_UP BL_DN[116] BL_DN[117]
+ BL_DN[118] BL_DN[119] BL_UP[116] BL_UP[117] BL_UP[118] BL_UP[119] GBL[29]
+ GBLB[29] GW[29] GWB[29] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_30 BLB_DN[120] BLB_DN[121] BLB_DN[122] BLB_DN[123] BLB_UP[120]
+ BLB_UP[121] BLB_UP[122] BLB_UP[123] BLEQ_DN BLEQ_UP BL_DN[120] BL_DN[121]
+ BL_DN[122] BL_DN[123] BL_UP[120] BL_UP[121] BL_UP[122] BL_UP[123] GBL[30]
+ GBLB[30] GW[30] GWB[30] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_31 BLB_DN[124] BLB_DN[125] BLB_DN[126] BLB_DN[127] BLB_UP[124]
+ BLB_UP[125] BLB_UP[126] BLB_UP[127] BLEQ_DN BLEQ_UP BL_DN[124] BL_DN[125]
+ BL_DN[126] BL_DN[127] BL_UP[124] BL_UP[125] BL_UP[126] BL_UP[127] GBL[31]
+ GBLB[31] GW[31] GWB[31] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_32 BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131] BLB_UP[128]
+ BLB_UP[129] BLB_UP[130] BLB_UP[131] BLEQ_DN BLEQ_UP BL_DN[128] BL_DN[129]
+ BL_DN[130] BL_DN[131] BL_UP[128] BL_UP[129] BL_UP[130] BL_UP[131] GBL[32]
+ GBLB[32] GW[32] GWB[32] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_33 BLB_DN[132] BLB_DN[133] BLB_DN[134] BLB_DN[135] BLB_UP[132]
+ BLB_UP[133] BLB_UP[134] BLB_UP[135] BLEQ_DN BLEQ_UP BL_DN[132] BL_DN[133]
+ BL_DN[134] BL_DN[135] BL_UP[132] BL_UP[133] BL_UP[134] BL_UP[135] GBL[33]
+ GBLB[33] GW[33] GWB[33] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_34 BLB_DN[136] BLB_DN[137] BLB_DN[138] BLB_DN[139] BLB_UP[136]
+ BLB_UP[137] BLB_UP[138] BLB_UP[139] BLEQ_DN BLEQ_UP BL_DN[136] BL_DN[137]
+ BL_DN[138] BL_DN[139] BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] GBL[34]
+ GBLB[34] GW[34] GWB[34] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_35 BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143] BLB_UP[140]
+ BLB_UP[141] BLB_UP[142] BLB_UP[143] BLEQ_DN BLEQ_UP BL_DN[140] BL_DN[141]
+ BL_DN[142] BL_DN[143] BL_UP[140] BL_UP[141] BL_UP[142] BL_UP[143] GBL[35]
+ GBLB[35] GW[35] GWB[35] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_36 BLB_DN[144] BLB_DN[145] BLB_DN[146] BLB_DN[147] BLB_UP[144]
+ BLB_UP[145] BLB_UP[146] BLB_UP[147] BLEQ_DN BLEQ_UP BL_DN[144] BL_DN[145]
+ BL_DN[146] BL_DN[147] BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147] GBL[36]
+ GBLB[36] GW[36] GWB[36] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_37 BLB_DN[148] BLB_DN[149] BLB_DN[150] BLB_DN[151] BLB_UP[148]
+ BLB_UP[149] BLB_UP[150] BLB_UP[151] BLEQ_DN BLEQ_UP BL_DN[148] BL_DN[149]
+ BL_DN[150] BL_DN[151] BL_UP[148] BL_UP[149] BL_UP[150] BL_UP[151] GBL[37]
+ GBLB[37] GW[37] GWB[37] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_38 BLB_DN[152] BLB_DN[153] BLB_DN[154] BLB_DN[155] BLB_UP[152]
+ BLB_UP[153] BLB_UP[154] BLB_UP[155] BLEQ_DN BLEQ_UP BL_DN[152] BL_DN[153]
+ BL_DN[154] BL_DN[155] BL_UP[152] BL_UP[153] BL_UP[154] BL_UP[155] GBL[38]
+ GBLB[38] GW[38] GWB[38] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_39 BLB_DN[156] BLB_DN[157] BLB_DN[158] BLB_DN[159] BLB_UP[156]
+ BLB_UP[157] BLB_UP[158] BLB_UP[159] BLEQ_DN BLEQ_UP BL_DN[156] BL_DN[157]
+ BL_DN[158] BL_DN[159] BL_UP[156] BL_UP[157] BL_UP[158] BL_UP[159] GBL[39]
+ GBLB[39] GW[39] GWB[39] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_40 BLB_DN[160] BLB_DN[161] BLB_DN[162] BLB_DN[163] BLB_UP[160]
+ BLB_UP[161] BLB_UP[162] BLB_UP[163] BLEQ_DN BLEQ_UP BL_DN[160] BL_DN[161]
+ BL_DN[162] BL_DN[163] BL_UP[160] BL_UP[161] BL_UP[162] BL_UP[163] GBL[40]
+ GBLB[40] GW[40] GWB[40] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_41 BLB_DN[164] BLB_DN[165] BLB_DN[166] BLB_DN[167] BLB_UP[164]
+ BLB_UP[165] BLB_UP[166] BLB_UP[167] BLEQ_DN BLEQ_UP BL_DN[164] BL_DN[165]
+ BL_DN[166] BL_DN[167] BL_UP[164] BL_UP[165] BL_UP[166] BL_UP[167] GBL[41]
+ GBLB[41] GW[41] GWB[41] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_42 BLB_DN[168] BLB_DN[169] BLB_DN[170] BLB_DN[171] BLB_UP[168]
+ BLB_UP[169] BLB_UP[170] BLB_UP[171] BLEQ_DN BLEQ_UP BL_DN[168] BL_DN[169]
+ BL_DN[170] BL_DN[171] BL_UP[168] BL_UP[169] BL_UP[170] BL_UP[171] GBL[42]
+ GBLB[42] GW[42] GWB[42] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_43 BLB_DN[172] BLB_DN[173] BLB_DN[174] BLB_DN[175] BLB_UP[172]
+ BLB_UP[173] BLB_UP[174] BLB_UP[175] BLEQ_DN BLEQ_UP BL_DN[172] BL_DN[173]
+ BL_DN[174] BL_DN[175] BL_UP[172] BL_UP[173] BL_UP[174] BL_UP[175] GBL[43]
+ GBLB[43] GW[43] GWB[43] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_44 BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179] BLB_UP[176]
+ BLB_UP[177] BLB_UP[178] BLB_UP[179] BLEQ_DN BLEQ_UP BL_DN[176] BL_DN[177]
+ BL_DN[178] BL_DN[179] BL_UP[176] BL_UP[177] BL_UP[178] BL_UP[179] GBL[44]
+ GBLB[44] GW[44] GWB[44] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_45 BLB_DN[180] BLB_DN[181] BLB_DN[182] BLB_DN[183] BLB_UP[180]
+ BLB_UP[181] BLB_UP[182] BLB_UP[183] BLEQ_DN BLEQ_UP BL_DN[180] BL_DN[181]
+ BL_DN[182] BL_DN[183] BL_UP[180] BL_UP[181] BL_UP[182] BL_UP[183] GBL[45]
+ GBLB[45] GW[45] GWB[45] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_46 BLB_DN[184] BLB_DN[185] BLB_DN[186] BLB_DN[187] BLB_UP[184]
+ BLB_UP[185] BLB_UP[186] BLB_UP[187] BLEQ_DN BLEQ_UP BL_DN[184] BL_DN[185]
+ BL_DN[186] BL_DN[187] BL_UP[184] BL_UP[185] BL_UP[186] BL_UP[187] GBL[46]
+ GBLB[46] GW[46] GWB[46] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_47 BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191] BLB_UP[188]
+ BLB_UP[189] BLB_UP[190] BLB_UP[191] BLEQ_DN BLEQ_UP BL_DN[188] BL_DN[189]
+ BL_DN[190] BL_DN[191] BL_UP[188] BL_UP[189] BL_UP[190] BL_UP[191] GBL[47]
+ GBLB[47] GW[47] GWB[47] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_48 BLB_DN[192] BLB_DN[193] BLB_DN[194] BLB_DN[195] BLB_UP[192]
+ BLB_UP[193] BLB_UP[194] BLB_UP[195] BLEQ_DN BLEQ_UP BL_DN[192] BL_DN[193]
+ BL_DN[194] BL_DN[195] BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] GBL[48]
+ GBLB[48] GW[48] GWB[48] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_49 BLB_DN[196] BLB_DN[197] BLB_DN[198] BLB_DN[199] BLB_UP[196]
+ BLB_UP[197] BLB_UP[198] BLB_UP[199] BLEQ_DN BLEQ_UP BL_DN[196] BL_DN[197]
+ BL_DN[198] BL_DN[199] BL_UP[196] BL_UP[197] BL_UP[198] BL_UP[199] GBL[49]
+ GBLB[49] GW[49] GWB[49] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_50 BLB_DN[200] BLB_DN[201] BLB_DN[202] BLB_DN[203] BLB_UP[200]
+ BLB_UP[201] BLB_UP[202] BLB_UP[203] BLEQ_DN BLEQ_UP BL_DN[200] BL_DN[201]
+ BL_DN[202] BL_DN[203] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203] GBL[50]
+ GBLB[50] GW[50] GWB[50] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_51 BLB_DN[204] BLB_DN[205] BLB_DN[206] BLB_DN[207] BLB_UP[204]
+ BLB_UP[205] BLB_UP[206] BLB_UP[207] BLEQ_DN BLEQ_UP BL_DN[204] BL_DN[205]
+ BL_DN[206] BL_DN[207] BL_UP[204] BL_UP[205] BL_UP[206] BL_UP[207] GBL[51]
+ GBLB[51] GW[51] GWB[51] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_52 BLB_DN[208] BLB_DN[209] BLB_DN[210] BLB_DN[211] BLB_UP[208]
+ BLB_UP[209] BLB_UP[210] BLB_UP[211] BLEQ_DN BLEQ_UP BL_DN[208] BL_DN[209]
+ BL_DN[210] BL_DN[211] BL_UP[208] BL_UP[209] BL_UP[210] BL_UP[211] GBL[52]
+ GBLB[52] GW[52] GWB[52] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_53 BLB_DN[212] BLB_DN[213] BLB_DN[214] BLB_DN[215] BLB_UP[212]
+ BLB_UP[213] BLB_UP[214] BLB_UP[215] BLEQ_DN BLEQ_UP BL_DN[212] BL_DN[213]
+ BL_DN[214] BL_DN[215] BL_UP[212] BL_UP[213] BL_UP[214] BL_UP[215] GBL[53]
+ GBLB[53] GW[53] GWB[53] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_54 BLB_DN[216] BLB_DN[217] BLB_DN[218] BLB_DN[219] BLB_UP[216]
+ BLB_UP[217] BLB_UP[218] BLB_UP[219] BLEQ_DN BLEQ_UP BL_DN[216] BL_DN[217]
+ BL_DN[218] BL_DN[219] BL_UP[216] BL_UP[217] BL_UP[218] BL_UP[219] GBL[54]
+ GBLB[54] GW[54] GWB[54] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_55 BLB_DN[220] BLB_DN[221] BLB_DN[222] BLB_DN[223] BLB_UP[220]
+ BLB_UP[221] BLB_UP[222] BLB_UP[223] BLEQ_DN BLEQ_UP BL_DN[220] BL_DN[221]
+ BL_DN[222] BL_DN[223] BL_UP[220] BL_UP[221] BL_UP[222] BL_UP[223] GBL[55]
+ GBLB[55] GW[55] GWB[55] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_56 BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227] BLB_UP[224]
+ BLB_UP[225] BLB_UP[226] BLB_UP[227] BLEQ_DN BLEQ_UP BL_DN[224] BL_DN[225]
+ BL_DN[226] BL_DN[227] BL_UP[224] BL_UP[225] BL_UP[226] BL_UP[227] GBL[56]
+ GBLB[56] GW[56] GWB[56] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_57 BLB_DN[228] BLB_DN[229] BLB_DN[230] BLB_DN[231] BLB_UP[228]
+ BLB_UP[229] BLB_UP[230] BLB_UP[231] BLEQ_DN BLEQ_UP BL_DN[228] BL_DN[229]
+ BL_DN[230] BL_DN[231] BL_UP[228] BL_UP[229] BL_UP[230] BL_UP[231] GBL[57]
+ GBLB[57] GW[57] GWB[57] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_58 BLB_DN[232] BLB_DN[233] BLB_DN[234] BLB_DN[235] BLB_UP[232]
+ BLB_UP[233] BLB_UP[234] BLB_UP[235] BLEQ_DN BLEQ_UP BL_DN[232] BL_DN[233]
+ BL_DN[234] BL_DN[235] BL_UP[232] BL_UP[233] BL_UP[234] BL_UP[235] GBL[58]
+ GBLB[58] GW[58] GWB[58] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_59 BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239] BLB_UP[236]
+ BLB_UP[237] BLB_UP[238] BLB_UP[239] BLEQ_DN BLEQ_UP BL_DN[236] BL_DN[237]
+ BL_DN[238] BL_DN[239] BL_UP[236] BL_UP[237] BL_UP[238] BL_UP[239] GBL[59]
+ GBLB[59] GW[59] GWB[59] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_60 BLB_DN[240] BLB_DN[241] BLB_DN[242] BLB_DN[243] BLB_UP[240]
+ BLB_UP[241] BLB_UP[242] BLB_UP[243] BLEQ_DN BLEQ_UP BL_DN[240] BL_DN[241]
+ BL_DN[242] BL_DN[243] BL_UP[240] BL_UP[241] BL_UP[242] BL_UP[243] GBL[60]
+ GBLB[60] GW[60] GWB[60] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_61 BLB_DN[244] BLB_DN[245] BLB_DN[246] BLB_DN[247] BLB_UP[244]
+ BLB_UP[245] BLB_UP[246] BLB_UP[247] BLEQ_DN BLEQ_UP BL_DN[244] BL_DN[245]
+ BL_DN[246] BL_DN[247] BL_UP[244] BL_UP[245] BL_UP[246] BL_UP[247] GBL[61]
+ GBLB[61] GW[61] GWB[61] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_62 BLB_DN[248] BLB_DN[249] BLB_DN[250] BLB_DN[251] BLB_UP[248]
+ BLB_UP[249] BLB_UP[250] BLB_UP[251] BLEQ_DN BLEQ_UP BL_DN[248] BL_DN[249]
+ BL_DN[250] BL_DN[251] BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] GBL[62]
+ GBLB[62] GW[62] GWB[62] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_63 BLB_DN[252] BLB_DN[253] BLB_DN[254] BLB_DN[255] BLB_UP[252]
+ BLB_UP[253] BLB_UP[254] BLB_UP[255] BLEQ_DN BLEQ_UP BL_DN[252] BL_DN[253]
+ BL_DN[254] BL_DN[255] BL_UP[252] BL_UP[253] BL_UP[254] BL_UP[255] GBL[63]
+ GBLB[63] GW[63] GWB[63] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_64 BLB_DN[256] BLB_DN[257] BLB_DN[258] BLB_DN[259] BLB_UP[256]
+ BLB_UP[257] BLB_UP[258] BLB_UP[259] BLEQ_DN BLEQ_UP BL_DN[256] BL_DN[257]
+ BL_DN[258] BL_DN[259] BL_UP[256] BL_UP[257] BL_UP[258] BL_UP[259] GBL[64]
+ GBLB[64] GW[64] GWB[64] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_65 BLB_DN[260] BLB_DN[261] BLB_DN[262] BLB_DN[263] BLB_UP[260]
+ BLB_UP[261] BLB_UP[262] BLB_UP[263] BLEQ_DN BLEQ_UP BL_DN[260] BL_DN[261]
+ BL_DN[262] BL_DN[263] BL_UP[260] BL_UP[261] BL_UP[262] BL_UP[263] GBL[65]
+ GBLB[65] GW[65] GWB[65] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_66 BLB_DN[264] BLB_DN[265] BLB_DN[266] BLB_DN[267] BLB_UP[264]
+ BLB_UP[265] BLB_UP[266] BLB_UP[267] BLEQ_DN BLEQ_UP BL_DN[264] BL_DN[265]
+ BL_DN[266] BL_DN[267] BL_UP[264] BL_UP[265] BL_UP[266] BL_UP[267] GBL[66]
+ GBLB[66] GW[66] GWB[66] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_67 BLB_DN[268] BLB_DN[269] BLB_DN[270] BLB_DN[271] BLB_UP[268]
+ BLB_UP[269] BLB_UP[270] BLB_UP[271] BLEQ_DN BLEQ_UP BL_DN[268] BL_DN[269]
+ BL_DN[270] BL_DN[271] BL_UP[268] BL_UP[269] BL_UP[270] BL_UP[271] GBL[67]
+ GBLB[67] GW[67] GWB[67] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_68 BLB_DN[272] BLB_DN[273] BLB_DN[274] BLB_DN[275] BLB_UP[272]
+ BLB_UP[273] BLB_UP[274] BLB_UP[275] BLEQ_DN BLEQ_UP BL_DN[272] BL_DN[273]
+ BL_DN[274] BL_DN[275] BL_UP[272] BL_UP[273] BL_UP[274] BL_UP[275] GBL[68]
+ GBLB[68] GW[68] GWB[68] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_69 BLB_DN[276] BLB_DN[277] BLB_DN[278] BLB_DN[279] BLB_UP[276]
+ BLB_UP[277] BLB_UP[278] BLB_UP[279] BLEQ_DN BLEQ_UP BL_DN[276] BL_DN[277]
+ BL_DN[278] BL_DN[279] BL_UP[276] BL_UP[277] BL_UP[278] BL_UP[279] GBL[69]
+ GBLB[69] GW[69] GWB[69] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_70 BLB_DN[280] BLB_DN[281] BLB_DN[282] BLB_DN[283] BLB_UP[280]
+ BLB_UP[281] BLB_UP[282] BLB_UP[283] BLEQ_DN BLEQ_UP BL_DN[280] BL_DN[281]
+ BL_DN[282] BL_DN[283] BL_UP[280] BL_UP[281] BL_UP[282] BL_UP[283] GBL[70]
+ GBLB[70] GW[70] GWB[70] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_71 BLB_DN[284] BLB_DN[285] BLB_DN[286] BLB_DN[287] BLB_UP[284]
+ BLB_UP[285] BLB_UP[286] BLB_UP[287] BLEQ_DN BLEQ_UP BL_DN[284] BL_DN[285]
+ BL_DN[286] BL_DN[287] BL_UP[284] BL_UP[285] BL_UP[286] BL_UP[287] GBL[71]
+ GBLB[71] GW[71] GWB[71] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_72 BLB_DN[288] BLB_DN[289] BLB_DN[290] BLB_DN[291] BLB_UP[288]
+ BLB_UP[289] BLB_UP[290] BLB_UP[291] BLEQ_DN BLEQ_UP BL_DN[288] BL_DN[289]
+ BL_DN[290] BL_DN[291] BL_UP[288] BL_UP[289] BL_UP[290] BL_UP[291] GBL[72]
+ GBLB[72] GW[72] GWB[72] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_73 BLB_DN[292] BLB_DN[293] BLB_DN[294] BLB_DN[295] BLB_UP[292]
+ BLB_UP[293] BLB_UP[294] BLB_UP[295] BLEQ_DN BLEQ_UP BL_DN[292] BL_DN[293]
+ BL_DN[294] BL_DN[295] BL_UP[292] BL_UP[293] BL_UP[294] BL_UP[295] GBL[73]
+ GBLB[73] GW[73] GWB[73] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_74 BLB_DN[296] BLB_DN[297] BLB_DN[298] BLB_DN[299] BLB_UP[296]
+ BLB_UP[297] BLB_UP[298] BLB_UP[299] BLEQ_DN BLEQ_UP BL_DN[296] BL_DN[297]
+ BL_DN[298] BL_DN[299] BL_UP[296] BL_UP[297] BL_UP[298] BL_UP[299] GBL[74]
+ GBLB[74] GW[74] GWB[74] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_75 BLB_DN[300] BLB_DN[301] BLB_DN[302] BLB_DN[303] BLB_UP[300]
+ BLB_UP[301] BLB_UP[302] BLB_UP[303] BLEQ_DN BLEQ_UP BL_DN[300] BL_DN[301]
+ BL_DN[302] BL_DN[303] BL_UP[300] BL_UP[301] BL_UP[302] BL_UP[303] GBL[75]
+ GBLB[75] GW[75] GWB[75] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_76 BLB_DN[304] BLB_DN[305] BLB_DN[306] BLB_DN[307] BLB_UP[304]
+ BLB_UP[305] BLB_UP[306] BLB_UP[307] BLEQ_DN BLEQ_UP BL_DN[304] BL_DN[305]
+ BL_DN[306] BL_DN[307] BL_UP[304] BL_UP[305] BL_UP[306] BL_UP[307] GBL[76]
+ GBLB[76] GW[76] GWB[76] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_77 BLB_DN[308] BLB_DN[309] BLB_DN[310] BLB_DN[311] BLB_UP[308]
+ BLB_UP[309] BLB_UP[310] BLB_UP[311] BLEQ_DN BLEQ_UP BL_DN[308] BL_DN[309]
+ BL_DN[310] BL_DN[311] BL_UP[308] BL_UP[309] BL_UP[310] BL_UP[311] GBL[77]
+ GBLB[77] GW[77] GWB[77] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_78 BLB_DN[312] BLB_DN[313] BLB_DN[314] BLB_DN[315] BLB_UP[312]
+ BLB_UP[313] BLB_UP[314] BLB_UP[315] BLEQ_DN BLEQ_UP BL_DN[312] BL_DN[313]
+ BL_DN[314] BL_DN[315] BL_UP[312] BL_UP[313] BL_UP[314] BL_UP[315] GBL[78]
+ GBLB[78] GW[78] GWB[78] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_79 BLB_DN[316] BLB_DN[317] BLB_DN[318] BLB_DN[319] BLB_UP[316]
+ BLB_UP[317] BLB_UP[318] BLB_UP[319] BLEQ_DN BLEQ_UP BL_DN[316] BL_DN[317]
+ BL_DN[318] BL_DN[319] BL_UP[316] BL_UP[317] BL_UP[318] BL_UP[319] GBL[79]
+ GBLB[79] GW[79] GWB[79] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_80 BLB_DN[320] BLB_DN[321] BLB_DN[322] BLB_DN[323] BLB_UP[320]
+ BLB_UP[321] BLB_UP[322] BLB_UP[323] BLEQ_DN BLEQ_UP BL_DN[320] BL_DN[321]
+ BL_DN[322] BL_DN[323] BL_UP[320] BL_UP[321] BL_UP[322] BL_UP[323] GBL[80]
+ GBLB[80] GW[80] GWB[80] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_81 BLB_DN[324] BLB_DN[325] BLB_DN[326] BLB_DN[327] BLB_UP[324]
+ BLB_UP[325] BLB_UP[326] BLB_UP[327] BLEQ_DN BLEQ_UP BL_DN[324] BL_DN[325]
+ BL_DN[326] BL_DN[327] BL_UP[324] BL_UP[325] BL_UP[326] BL_UP[327] GBL[81]
+ GBLB[81] GW[81] GWB[81] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_82 BLB_DN[328] BLB_DN[329] BLB_DN[330] BLB_DN[331] BLB_UP[328]
+ BLB_UP[329] BLB_UP[330] BLB_UP[331] BLEQ_DN BLEQ_UP BL_DN[328] BL_DN[329]
+ BL_DN[330] BL_DN[331] BL_UP[328] BL_UP[329] BL_UP[330] BL_UP[331] GBL[82]
+ GBLB[82] GW[82] GWB[82] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_83 BLB_DN[332] BLB_DN[333] BLB_DN[334] BLB_DN[335] BLB_UP[332]
+ BLB_UP[333] BLB_UP[334] BLB_UP[335] BLEQ_DN BLEQ_UP BL_DN[332] BL_DN[333]
+ BL_DN[334] BL_DN[335] BL_UP[332] BL_UP[333] BL_UP[334] BL_UP[335] GBL[83]
+ GBLB[83] GW[83] GWB[83] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_84 BLB_DN[336] BLB_DN[337] BLB_DN[338] BLB_DN[339] BLB_UP[336]
+ BLB_UP[337] BLB_UP[338] BLB_UP[339] BLEQ_DN BLEQ_UP BL_DN[336] BL_DN[337]
+ BL_DN[338] BL_DN[339] BL_UP[336] BL_UP[337] BL_UP[338] BL_UP[339] GBL[84]
+ GBLB[84] GW[84] GWB[84] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_85 BLB_DN[340] BLB_DN[341] BLB_DN[342] BLB_DN[343] BLB_UP[340]
+ BLB_UP[341] BLB_UP[342] BLB_UP[343] BLEQ_DN BLEQ_UP BL_DN[340] BL_DN[341]
+ BL_DN[342] BL_DN[343] BL_UP[340] BL_UP[341] BL_UP[342] BL_UP[343] GBL[85]
+ GBLB[85] GW[85] GWB[85] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_86 BLB_DN[344] BLB_DN[345] BLB_DN[346] BLB_DN[347] BLB_UP[344]
+ BLB_UP[345] BLB_UP[346] BLB_UP[347] BLEQ_DN BLEQ_UP BL_DN[344] BL_DN[345]
+ BL_DN[346] BL_DN[347] BL_UP[344] BL_UP[345] BL_UP[346] BL_UP[347] GBL[86]
+ GBLB[86] GW[86] GWB[86] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_87 BLB_DN[348] BLB_DN[349] BLB_DN[350] BLB_DN[351] BLB_UP[348]
+ BLB_UP[349] BLB_UP[350] BLB_UP[351] BLEQ_DN BLEQ_UP BL_DN[348] BL_DN[349]
+ BL_DN[350] BL_DN[351] BL_UP[348] BL_UP[349] BL_UP[350] BL_UP[351] GBL[87]
+ GBLB[87] GW[87] GWB[87] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_88 BLB_DN[352] BLB_DN[353] BLB_DN[354] BLB_DN[355] BLB_UP[352]
+ BLB_UP[353] BLB_UP[354] BLB_UP[355] BLEQ_DN BLEQ_UP BL_DN[352] BL_DN[353]
+ BL_DN[354] BL_DN[355] BL_UP[352] BL_UP[353] BL_UP[354] BL_UP[355] GBL[88]
+ GBLB[88] GW[88] GWB[88] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_89 BLB_DN[356] BLB_DN[357] BLB_DN[358] BLB_DN[359] BLB_UP[356]
+ BLB_UP[357] BLB_UP[358] BLB_UP[359] BLEQ_DN BLEQ_UP BL_DN[356] BL_DN[357]
+ BL_DN[358] BL_DN[359] BL_UP[356] BL_UP[357] BL_UP[358] BL_UP[359] GBL[89]
+ GBLB[89] GW[89] GWB[89] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_90 BLB_DN[360] BLB_DN[361] BLB_DN[362] BLB_DN[363] BLB_UP[360]
+ BLB_UP[361] BLB_UP[362] BLB_UP[363] BLEQ_DN BLEQ_UP BL_DN[360] BL_DN[361]
+ BL_DN[362] BL_DN[363] BL_UP[360] BL_UP[361] BL_UP[362] BL_UP[363] GBL[90]
+ GBLB[90] GW[90] GWB[90] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_91 BLB_DN[364] BLB_DN[365] BLB_DN[366] BLB_DN[367] BLB_UP[364]
+ BLB_UP[365] BLB_UP[366] BLB_UP[367] BLEQ_DN BLEQ_UP BL_DN[364] BL_DN[365]
+ BL_DN[366] BL_DN[367] BL_UP[364] BL_UP[365] BL_UP[366] BL_UP[367] GBL[91]
+ GBLB[91] GW[91] GWB[91] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_92 BLB_DN[368] BLB_DN[369] BLB_DN[370] BLB_DN[371] BLB_UP[368]
+ BLB_UP[369] BLB_UP[370] BLB_UP[371] BLEQ_DN BLEQ_UP BL_DN[368] BL_DN[369]
+ BL_DN[370] BL_DN[371] BL_UP[368] BL_UP[369] BL_UP[370] BL_UP[371] GBL[92]
+ GBLB[92] GW[92] GWB[92] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_93 BLB_DN[372] BLB_DN[373] BLB_DN[374] BLB_DN[375] BLB_UP[372]
+ BLB_UP[373] BLB_UP[374] BLB_UP[375] BLEQ_DN BLEQ_UP BL_DN[372] BL_DN[373]
+ BL_DN[374] BL_DN[375] BL_UP[372] BL_UP[373] BL_UP[374] BL_UP[375] GBL[93]
+ GBLB[93] GW[93] GWB[93] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_94 BLB_DN[376] BLB_DN[377] BLB_DN[378] BLB_DN[379] BLB_UP[376]
+ BLB_UP[377] BLB_UP[378] BLB_UP[379] BLEQ_DN BLEQ_UP BL_DN[376] BL_DN[377]
+ BL_DN[378] BL_DN[379] BL_UP[376] BL_UP[377] BL_UP[378] BL_UP[379] GBL[94]
+ GBLB[94] GW[94] GWB[94] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_95 BLB_DN[380] BLB_DN[381] BLB_DN[382] BLB_DN[383] BLB_UP[380]
+ BLB_UP[381] BLB_UP[382] BLB_UP[383] BLEQ_DN BLEQ_UP BL_DN[380] BL_DN[381]
+ BL_DN[382] BL_DN[383] BL_UP[380] BL_UP[381] BL_UP[382] BL_UP[383] GBL[95]
+ GBLB[95] GW[95] GWB[95] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_96 BLB_DN[384] BLB_DN[385] BLB_DN[386] BLB_DN[387] BLB_UP[384]
+ BLB_UP[385] BLB_UP[386] BLB_UP[387] BLEQ_DN BLEQ_UP BL_DN[384] BL_DN[385]
+ BL_DN[386] BL_DN[387] BL_UP[384] BL_UP[385] BL_UP[386] BL_UP[387] GBL[96]
+ GBLB[96] GW[96] GWB[96] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_97 BLB_DN[388] BLB_DN[389] BLB_DN[390] BLB_DN[391] BLB_UP[388]
+ BLB_UP[389] BLB_UP[390] BLB_UP[391] BLEQ_DN BLEQ_UP BL_DN[388] BL_DN[389]
+ BL_DN[390] BL_DN[391] BL_UP[388] BL_UP[389] BL_UP[390] BL_UP[391] GBL[97]
+ GBLB[97] GW[97] GWB[97] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_98 BLB_DN[392] BLB_DN[393] BLB_DN[394] BLB_DN[395] BLB_UP[392]
+ BLB_UP[393] BLB_UP[394] BLB_UP[395] BLEQ_DN BLEQ_UP BL_DN[392] BL_DN[393]
+ BL_DN[394] BL_DN[395] BL_UP[392] BL_UP[393] BL_UP[394] BL_UP[395] GBL[98]
+ GBLB[98] GW[98] GWB[98] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_99 BLB_DN[396] BLB_DN[397] BLB_DN[398] BLB_DN[399] BLB_UP[396]
+ BLB_UP[397] BLB_UP[398] BLB_UP[399] BLEQ_DN BLEQ_UP BL_DN[396] BL_DN[397]
+ BL_DN[398] BL_DN[399] BL_UP[396] BL_UP[397] BL_UP[398] BL_UP[399] GBL[99]
+ GBLB[99] GW[99] GWB[99] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_100 BLB_DN[400] BLB_DN[401] BLB_DN[402] BLB_DN[403] BLB_UP[400]
+ BLB_UP[401] BLB_UP[402] BLB_UP[403] BLEQ_DN BLEQ_UP BL_DN[400] BL_DN[401]
+ BL_DN[402] BL_DN[403] BL_UP[400] BL_UP[401] BL_UP[402] BL_UP[403] GBL[100]
+ GBLB[100] GW[100] GWB[100] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_101 BLB_DN[404] BLB_DN[405] BLB_DN[406] BLB_DN[407] BLB_UP[404]
+ BLB_UP[405] BLB_UP[406] BLB_UP[407] BLEQ_DN BLEQ_UP BL_DN[404] BL_DN[405]
+ BL_DN[406] BL_DN[407] BL_UP[404] BL_UP[405] BL_UP[406] BL_UP[407] GBL[101]
+ GBLB[101] GW[101] GWB[101] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_102 BLB_DN[408] BLB_DN[409] BLB_DN[410] BLB_DN[411] BLB_UP[408]
+ BLB_UP[409] BLB_UP[410] BLB_UP[411] BLEQ_DN BLEQ_UP BL_DN[408] BL_DN[409]
+ BL_DN[410] BL_DN[411] BL_UP[408] BL_UP[409] BL_UP[410] BL_UP[411] GBL[102]
+ GBLB[102] GW[102] GWB[102] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_103 BLB_DN[412] BLB_DN[413] BLB_DN[414] BLB_DN[415] BLB_UP[412]
+ BLB_UP[413] BLB_UP[414] BLB_UP[415] BLEQ_DN BLEQ_UP BL_DN[412] BL_DN[413]
+ BL_DN[414] BL_DN[415] BL_UP[412] BL_UP[413] BL_UP[414] BL_UP[415] GBL[103]
+ GBLB[103] GW[103] GWB[103] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_104 BLB_DN[416] BLB_DN[417] BLB_DN[418] BLB_DN[419] BLB_UP[416]
+ BLB_UP[417] BLB_UP[418] BLB_UP[419] BLEQ_DN BLEQ_UP BL_DN[416] BL_DN[417]
+ BL_DN[418] BL_DN[419] BL_UP[416] BL_UP[417] BL_UP[418] BL_UP[419] GBL[104]
+ GBLB[104] GW[104] GWB[104] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_105 BLB_DN[420] BLB_DN[421] BLB_DN[422] BLB_DN[423] BLB_UP[420]
+ BLB_UP[421] BLB_UP[422] BLB_UP[423] BLEQ_DN BLEQ_UP BL_DN[420] BL_DN[421]
+ BL_DN[422] BL_DN[423] BL_UP[420] BL_UP[421] BL_UP[422] BL_UP[423] GBL[105]
+ GBLB[105] GW[105] GWB[105] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_106 BLB_DN[424] BLB_DN[425] BLB_DN[426] BLB_DN[427] BLB_UP[424]
+ BLB_UP[425] BLB_UP[426] BLB_UP[427] BLEQ_DN BLEQ_UP BL_DN[424] BL_DN[425]
+ BL_DN[426] BL_DN[427] BL_UP[424] BL_UP[425] BL_UP[426] BL_UP[427] GBL[106]
+ GBLB[106] GW[106] GWB[106] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_107 BLB_DN[428] BLB_DN[429] BLB_DN[430] BLB_DN[431] BLB_UP[428]
+ BLB_UP[429] BLB_UP[430] BLB_UP[431] BLEQ_DN BLEQ_UP BL_DN[428] BL_DN[429]
+ BL_DN[430] BL_DN[431] BL_UP[428] BL_UP[429] BL_UP[430] BL_UP[431] GBL[107]
+ GBLB[107] GW[107] GWB[107] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_108 BLB_DN[432] BLB_DN[433] BLB_DN[434] BLB_DN[435] BLB_UP[432]
+ BLB_UP[433] BLB_UP[434] BLB_UP[435] BLEQ_DN BLEQ_UP BL_DN[432] BL_DN[433]
+ BL_DN[434] BL_DN[435] BL_UP[432] BL_UP[433] BL_UP[434] BL_UP[435] GBL[108]
+ GBLB[108] GW[108] GWB[108] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_109 BLB_DN[436] BLB_DN[437] BLB_DN[438] BLB_DN[439] BLB_UP[436]
+ BLB_UP[437] BLB_UP[438] BLB_UP[439] BLEQ_DN BLEQ_UP BL_DN[436] BL_DN[437]
+ BL_DN[438] BL_DN[439] BL_UP[436] BL_UP[437] BL_UP[438] BL_UP[439] GBL[109]
+ GBLB[109] GW[109] GWB[109] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_110 BLB_DN[440] BLB_DN[441] BLB_DN[442] BLB_DN[443] BLB_UP[440]
+ BLB_UP[441] BLB_UP[442] BLB_UP[443] BLEQ_DN BLEQ_UP BL_DN[440] BL_DN[441]
+ BL_DN[442] BL_DN[443] BL_UP[440] BL_UP[441] BL_UP[442] BL_UP[443] GBL[110]
+ GBLB[110] GW[110] GWB[110] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_111 BLB_DN[444] BLB_DN[445] BLB_DN[446] BLB_DN[447] BLB_UP[444]
+ BLB_UP[445] BLB_UP[446] BLB_UP[447] BLEQ_DN BLEQ_UP BL_DN[444] BL_DN[445]
+ BL_DN[446] BL_DN[447] BL_UP[444] BL_UP[445] BL_UP[446] BL_UP[447] GBL[111]
+ GBLB[111] GW[111] GWB[111] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_112 BLB_DN[448] BLB_DN[449] BLB_DN[450] BLB_DN[451] BLB_UP[448]
+ BLB_UP[449] BLB_UP[450] BLB_UP[451] BLEQ_DN BLEQ_UP BL_DN[448] BL_DN[449]
+ BL_DN[450] BL_DN[451] BL_UP[448] BL_UP[449] BL_UP[450] BL_UP[451] GBL[112]
+ GBLB[112] GW[112] GWB[112] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_113 BLB_DN[452] BLB_DN[453] BLB_DN[454] BLB_DN[455] BLB_UP[452]
+ BLB_UP[453] BLB_UP[454] BLB_UP[455] BLEQ_DN BLEQ_UP BL_DN[452] BL_DN[453]
+ BL_DN[454] BL_DN[455] BL_UP[452] BL_UP[453] BL_UP[454] BL_UP[455] GBL[113]
+ GBLB[113] GW[113] GWB[113] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_114 BLB_DN[456] BLB_DN[457] BLB_DN[458] BLB_DN[459] BLB_UP[456]
+ BLB_UP[457] BLB_UP[458] BLB_UP[459] BLEQ_DN BLEQ_UP BL_DN[456] BL_DN[457]
+ BL_DN[458] BL_DN[459] BL_UP[456] BL_UP[457] BL_UP[458] BL_UP[459] GBL[114]
+ GBLB[114] GW[114] GWB[114] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_115 BLB_DN[460] BLB_DN[461] BLB_DN[462] BLB_DN[463] BLB_UP[460]
+ BLB_UP[461] BLB_UP[462] BLB_UP[463] BLEQ_DN BLEQ_UP BL_DN[460] BL_DN[461]
+ BL_DN[462] BL_DN[463] BL_UP[460] BL_UP[461] BL_UP[462] BL_UP[463] GBL[115]
+ GBLB[115] GW[115] GWB[115] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_116 BLB_DN[464] BLB_DN[465] BLB_DN[466] BLB_DN[467] BLB_UP[464]
+ BLB_UP[465] BLB_UP[466] BLB_UP[467] BLEQ_DN BLEQ_UP BL_DN[464] BL_DN[465]
+ BL_DN[466] BL_DN[467] BL_UP[464] BL_UP[465] BL_UP[466] BL_UP[467] GBL[116]
+ GBLB[116] GW[116] GWB[116] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_117 BLB_DN[468] BLB_DN[469] BLB_DN[470] BLB_DN[471] BLB_UP[468]
+ BLB_UP[469] BLB_UP[470] BLB_UP[471] BLEQ_DN BLEQ_UP BL_DN[468] BL_DN[469]
+ BL_DN[470] BL_DN[471] BL_UP[468] BL_UP[469] BL_UP[470] BL_UP[471] GBL[117]
+ GBLB[117] GW[117] GWB[117] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_118 BLB_DN[472] BLB_DN[473] BLB_DN[474] BLB_DN[475] BLB_UP[472]
+ BLB_UP[473] BLB_UP[474] BLB_UP[475] BLEQ_DN BLEQ_UP BL_DN[472] BL_DN[473]
+ BL_DN[474] BL_DN[475] BL_UP[472] BL_UP[473] BL_UP[474] BL_UP[475] GBL[118]
+ GBLB[118] GW[118] GWB[118] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_119 BLB_DN[476] BLB_DN[477] BLB_DN[478] BLB_DN[479] BLB_UP[476]
+ BLB_UP[477] BLB_UP[478] BLB_UP[479] BLEQ_DN BLEQ_UP BL_DN[476] BL_DN[477]
+ BL_DN[478] BL_DN[479] BL_UP[476] BL_UP[477] BL_UP[478] BL_UP[479] GBL[119]
+ GBLB[119] GW[119] GWB[119] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_120 BLB_DN[480] BLB_DN[481] BLB_DN[482] BLB_DN[483] BLB_UP[480]
+ BLB_UP[481] BLB_UP[482] BLB_UP[483] BLEQ_DN BLEQ_UP BL_DN[480] BL_DN[481]
+ BL_DN[482] BL_DN[483] BL_UP[480] BL_UP[481] BL_UP[482] BL_UP[483] GBL[120]
+ GBLB[120] GW[120] GWB[120] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_121 BLB_DN[484] BLB_DN[485] BLB_DN[486] BLB_DN[487] BLB_UP[484]
+ BLB_UP[485] BLB_UP[486] BLB_UP[487] BLEQ_DN BLEQ_UP BL_DN[484] BL_DN[485]
+ BL_DN[486] BL_DN[487] BL_UP[484] BL_UP[485] BL_UP[486] BL_UP[487] GBL[121]
+ GBLB[121] GW[121] GWB[121] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_122 BLB_DN[488] BLB_DN[489] BLB_DN[490] BLB_DN[491] BLB_UP[488]
+ BLB_UP[489] BLB_UP[490] BLB_UP[491] BLEQ_DN BLEQ_UP BL_DN[488] BL_DN[489]
+ BL_DN[490] BL_DN[491] BL_UP[488] BL_UP[489] BL_UP[490] BL_UP[491] GBL[122]
+ GBLB[122] GW[122] GWB[122] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_123 BLB_DN[492] BLB_DN[493] BLB_DN[494] BLB_DN[495] BLB_UP[492]
+ BLB_UP[493] BLB_UP[494] BLB_UP[495] BLEQ_DN BLEQ_UP BL_DN[492] BL_DN[493]
+ BL_DN[494] BL_DN[495] BL_UP[492] BL_UP[493] BL_UP[494] BL_UP[495] GBL[123]
+ GBLB[123] GW[123] GWB[123] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_124 BLB_DN[496] BLB_DN[497] BLB_DN[498] BLB_DN[499] BLB_UP[496]
+ BLB_UP[497] BLB_UP[498] BLB_UP[499] BLEQ_DN BLEQ_UP BL_DN[496] BL_DN[497]
+ BL_DN[498] BL_DN[499] BL_UP[496] BL_UP[497] BL_UP[498] BL_UP[499] GBL[124]
+ GBLB[124] GW[124] GWB[124] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_125 BLB_DN[500] BLB_DN[501] BLB_DN[502] BLB_DN[503] BLB_UP[500]
+ BLB_UP[501] BLB_UP[502] BLB_UP[503] BLEQ_DN BLEQ_UP BL_DN[500] BL_DN[501]
+ BL_DN[502] BL_DN[503] BL_UP[500] BL_UP[501] BL_UP[502] BL_UP[503] GBL[125]
+ GBLB[125] GW[125] GWB[125] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_126 BLB_DN[504] BLB_DN[505] BLB_DN[506] BLB_DN[507] BLB_UP[504]
+ BLB_UP[505] BLB_UP[506] BLB_UP[507] BLEQ_DN BLEQ_UP BL_DN[504] BL_DN[505]
+ BL_DN[506] BL_DN[507] BL_UP[504] BL_UP[505] BL_UP[506] BL_UP[507] GBL[126]
+ GBLB[126] GW[126] GWB[126] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
XLIO_M4_127 BLB_DN[508] BLB_DN[509] BLB_DN[510] BLB_DN[511] BLB_UP[508]
+ BLB_UP[509] BLB_UP[510] BLB_UP[511] BLEQ_DN BLEQ_UP BL_DN[508] BL_DN[509]
+ BL_DN[510] BL_DN[511] BL_UP[508] BL_UP[509] BL_UP[510] BL_UP[511] GBL[127]
+ GBLB[127] GW[127] GWB[127] PREBG SAEB VDDI VSSI Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] SDBM200W80_LIO_M4
.ENDS

.SUBCKT SDBM200W80_WL_TRK WL_TK BL_TK SLP_BUF TIEH TIEL VDDI VSSI
XTKWL_2X2_RL0 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL1 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL2 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL3 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL4 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL5 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL6 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL7 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL8 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL9 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL10 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL11 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL12 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL13 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL14 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL15 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL16 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL17 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL18 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL19 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL20 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL21 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL22 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL23 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL24 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL25 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL26 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL27 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL28 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL29 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL30 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL31 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL32 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL33 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL34 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL35 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL36 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL37 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL38 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL39 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL40 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL41 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL42 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL43 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL44 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL45 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL46 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL47 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL48 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL49 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL50 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL51 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL52 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL53 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL54 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL55 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL56 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL57 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_RL58 VDDI VSSI WL_TK WL_TK SDBM200W80_TKWL_2X2
XTKWL_2X2_ISO VDDI VSSI WL_TK WL_TK TIEL TIEL SDBM200W80_TKWL_2X2_ISO
XTKWL_2X2_RR0 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR1 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR2 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR3 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR4 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR5 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR6 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR7 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR8 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR9 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR10 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR11 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR12 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR13 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR14 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR15 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR16 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR17 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR18 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR19 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR20 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR21 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR22 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR23 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR24 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR25 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR26 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR27 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR28 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR29 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR30 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR31 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR32 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR33 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR34 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR35 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR36 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR37 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR38 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR39 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR40 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR41 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR42 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR43 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR44 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR45 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR46 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR47 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR48 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR49 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR50 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR51 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR52 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR53 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR54 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR55 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR56 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR57 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR58 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR59 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR60 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR61 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR62 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR63 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR64 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR65 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR66 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR67 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_RR68 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKBL_TRKPRE BL_TK WL_TK VDDI VSSI TIEH TIEL SDBM200W80_TKBL_TRKPRE
XTKWL_2X2_L0 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L1 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L2 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L3 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L4 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L5 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L6 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L7 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L8 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L9 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L10 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L11 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L12 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L13 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L14 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L15 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L16 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L17 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L18 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L19 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L20 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L21 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L22 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L23 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L24 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L25 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L26 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L27 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L28 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L29 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L30 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L31 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L32 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L33 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L34 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L35 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L36 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L37 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L38 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L39 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L40 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L41 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L42 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L43 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L44 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L45 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L46 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L47 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L48 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L49 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L50 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L51 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L52 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L53 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L54 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L55 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L56 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L57 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L58 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L59 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L60 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L61 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L62 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L63 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L64 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L65 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L66 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L67 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L68 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L69 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L70 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L71 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L72 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L73 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L74 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L75 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L76 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L77 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L78 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L79 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L80 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L81 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L82 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L83 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L84 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L85 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L86 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L87 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L88 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L89 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L90 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L91 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L92 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L93 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L94 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L95 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L96 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L97 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L98 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L99 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L100 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L101 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L102 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L103 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L104 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L105 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L106 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L107 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L108 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L109 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L110 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L111 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L112 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L113 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L114 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L115 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L116 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L117 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L118 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L119 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L120 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L121 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L122 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L123 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L124 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L125 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L126 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
XTKWL_2X2_L127 VDDI VSSI TIEL TIEL SDBM200W80_TKWL_2X2
.ENDS

.SUBCKT SDBM200W80_TRACKING WL_TK SLP_BUF BL_TK WL[0] WL[1] WL[2] WL[3] WL[4]
+ WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16]
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27]
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38]
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49]
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60]
+ WL[61] WL[62] WL[63] VDDI VSSI
XWL_TRK WL_TK BL_TK SLP_BUF TIEH TIEL VDDI VSSI SDBM200W80_WL_TRK
X0TRKNORX2_0 BL_TK VDDI VSSI WL[0] WL[1] WL_TK FLOAT1[0] NET[0] FLOAT3
+ NET_TRKBL[0] FLOAT5 TIEH SDBM200W80_TRKNORX2
X1TRKNORX2_1 BL_TK VDDI VSSI WL[2] WL[3] WL_TK FLOAT1[1] NET[1] NET[0]
+ NET_TRKBL[1] NET_TRKBL[0] TIEH SDBM200W80_TRKNORX2
X2TRKNORX2_2 BL_TK VDDI VSSI WL[4] WL[5] WL_TK FLOAT1[2] NET[2] NET[1]
+ NET_TRKBL[2] NET_TRKBL[1] TIEH SDBM200W80_TRKNORX2
X3TRKNORX2_3 BL_TK VDDI VSSI WL[6] WL[7] WL_TK FLOAT1[3] NET[3] NET[2]
+ NET_TRKBL[3] NET_TRKBL[2] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_4 BL_TK VDDI VSSI WL[8] WL[9] TIEL FLOAT1[4] NET[4] NET[3]
+ NET_TRKBL[4] NET_TRKBL[3] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_5 BL_TK VDDI VSSI WL[10] WL[11] TIEL FLOAT1[5] NET[5] NET[4]
+ NET_TRKBL[5] NET_TRKBL[4] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_6 BL_TK VDDI VSSI WL[12] WL[13] TIEL FLOAT1[6] NET[6] NET[5]
+ NET_TRKBL[6] NET_TRKBL[5] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_7 BL_TK VDDI VSSI WL[14] WL[15] TIEL FLOAT1[7] NET[7] NET[6]
+ NET_TRKBL[7] NET_TRKBL[6] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_8 BL_TK VDDI VSSI WL[16] WL[17] TIEL FLOAT1[8] NET[8] NET[7]
+ NET_TRKBL[8] NET_TRKBL[7] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_9 BL_TK VDDI VSSI WL[18] WL[19] TIEL FLOAT1[9] NET[9] NET[8]
+ NET_TRKBL[9] NET_TRKBL[8] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_10 BL_TK VDDI VSSI WL[20] WL[21] TIEL FLOAT1[10] NET[10] NET[9]
+ NET_TRKBL[10] NET_TRKBL[9] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_11 BL_TK VDDI VSSI WL[22] WL[23] TIEL FLOAT1[11] NET[11] NET[10]
+ NET_TRKBL[11] NET_TRKBL[10] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_12 BL_TK VDDI VSSI WL[24] WL[25] TIEL FLOAT1[12] NET[12] NET[11]
+ NET_TRKBL[12] NET_TRKBL[11] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_13 BL_TK VDDI VSSI WL[26] WL[27] TIEL FLOAT1[13] NET[13] NET[12]
+ NET_TRKBL[13] NET_TRKBL[12] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_14 BL_TK VDDI VSSI WL[28] WL[29] TIEL FLOAT1[14] NET[14] NET[13]
+ NET_TRKBL[14] NET_TRKBL[13] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_15 BL_TK VDDI VSSI WL[30] WL[31] TIEL FLOAT1[15] NET[15] NET[14]
+ NET_TRKBL[15] NET_TRKBL[14] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_16 BL_TK VDDI VSSI WL[32] WL[33] TIEL FLOAT1[16] NET[16] NET[15]
+ NET_TRKBL[16] NET_TRKBL[15] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_17 BL_TK VDDI VSSI WL[34] WL[35] TIEL FLOAT1[17] NET[17] NET[16]
+ NET_TRKBL[17] NET_TRKBL[16] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_18 BL_TK VDDI VSSI WL[36] WL[37] TIEL FLOAT1[18] NET[18] NET[17]
+ NET_TRKBL[18] NET_TRKBL[17] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_19 BL_TK VDDI VSSI WL[38] WL[39] TIEL FLOAT1[19] NET[19] NET[18]
+ NET_TRKBL[19] NET_TRKBL[18] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_20 BL_TK VDDI VSSI WL[40] WL[41] TIEL FLOAT1[20] NET[20] NET[19]
+ NET_TRKBL[20] NET_TRKBL[19] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_21 BL_TK VDDI VSSI WL[42] WL[43] TIEL FLOAT1[21] NET[21] NET[20]
+ NET_TRKBL[21] NET_TRKBL[20] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_22 BL_TK VDDI VSSI WL[44] WL[45] TIEL FLOAT1[22] NET[22] NET[21]
+ NET_TRKBL[22] NET_TRKBL[21] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_23 BL_TK VDDI VSSI WL[46] WL[47] TIEL FLOAT1[23] NET[23] NET[22]
+ NET_TRKBL[23] NET_TRKBL[22] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_24 BL_TK VDDI VSSI WL[48] WL[49] TIEL FLOAT1[24] NET[24] NET[23]
+ NET_TRKBL[24] NET_TRKBL[23] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_25 BL_TK VDDI VSSI WL[50] WL[51] TIEL FLOAT1[25] NET[25] NET[24]
+ NET_TRKBL[25] NET_TRKBL[24] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_26 BL_TK VDDI VSSI WL[52] WL[53] TIEL FLOAT1[26] NET[26] NET[25]
+ NET_TRKBL[26] NET_TRKBL[25] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_27 BL_TK VDDI VSSI WL[54] WL[55] TIEL FLOAT1[27] NET[27] NET[26]
+ NET_TRKBL[27] NET_TRKBL[26] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_28 BL_TK VDDI VSSI WL[56] WL[57] TIEL FLOAT1[28] NET[28] NET[27]
+ NET_TRKBL[28] NET_TRKBL[27] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_29 BL_TK VDDI VSSI WL[58] WL[59] TIEL FLOAT1[29] NET[29] NET[28]
+ NET_TRKBL[29] NET_TRKBL[28] TIEH SDBM200W80_TRKNORX2
X4TRKNORX2_30 BL_TK VDDI VSSI WL[60] WL[61] TIEL FLOAT1[30] NET[30] NET[29]
+ NET_TRKBL[30] NET_TRKBL[29] TIEH SDBM200W80_TRKNORX2
X5TRKNORX2_31 BL_TK VDDI VSSI WL[62] WL[63] TIEL FLOAT1[31] NET[31] NET[30]
+ NET_TRKBL[31] NET_TRKBL[30] TIEH SDBM200W80_TRKNORX2
.ENDS

.SUBCKT SDBM200W80_BANK_0_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6]
+ GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16]
+ GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25]
+ GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34]
+ GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43]
+ GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52]
+ GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61]
+ GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69] GBL[70]
+ GBL[71] GBL[72] GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78] GBL[79]
+ GBL[80] GBL[81] GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87] GBL[88]
+ GBL[89] GBL[90] GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96] GBL[97]
+ GBL[98] GBL[99] GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105] GBL[106]
+ GBL[107] GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113] GBL[114]
+ GBL[115] GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121] GBL[122]
+ GBL[123] GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2] GBLB[3]
+ GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12]
+ GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20]
+ GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28]
+ GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36]
+ GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44]
+ GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52]
+ GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60]
+ GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67] GBLB[68]
+ GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75] GBLB[76]
+ GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83] GBLB[84]
+ GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91] GBLB[92]
+ GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99] GBLB[100]
+ GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106] GBLB[107]
+ GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113] GBLB[114]
+ GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120] GBLB[121]
+ GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0] GW[1] GW[2]
+ GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14]
+ GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25]
+ GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36]
+ GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47]
+ GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58]
+ GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67] GW[68] GW[69]
+ GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78] GW[79] GW[80]
+ GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89] GW[90] GW[91]
+ GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100] GW[101]
+ GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109] GW[110]
+ GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118] GW[119]
+ GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65]
+ GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74]
+ GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83]
+ GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92]
+ GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101]
+ GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109]
+ GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117]
+ GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125]
+ GWB[126] GWB[127] SLP_LCTRL WLP_SAE DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1]
+ DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] BL_TK WL_TK VDDI VSSI WLP_SAE_TK
XTRACKING WL_TK SLP_LCTRL BL_TK WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7]
+ WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18]
+ WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29]
+ WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40]
+ WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51]
+ WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62]
+ WL[63] VDDI VSSI SDBM200W80_TRACKING
XLIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36]
+ GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45]
+ GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54]
+ GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63]
+ GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69] GBL[70] GBL[71] GBL[72]
+ GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78] GBL[79] GBL[80] GBL[81]
+ GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87] GBL[88] GBL[89] GBL[90]
+ GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96] GBL[97] GBL[98] GBL[99]
+ GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105] GBL[106] GBL[107]
+ GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113] GBL[114] GBL[115]
+ GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121] GBL[122] GBL[123]
+ GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37]
+ GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45]
+ GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53]
+ GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61]
+ GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67] GBLB[68] GBLB[69]
+ GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75] GBLB[76] GBLB[77]
+ GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83] GBLB[84] GBLB[85]
+ GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91] GBLB[92] GBLB[93]
+ GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99] GBLB[100] GBLB[101]
+ GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106] GBLB[107] GBLB[108]
+ GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113] GBLB[114] GBLB[115]
+ GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120] GBLB[121] GBLB[122]
+ GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] LIOPD WL[0] WL[1] WL[2]
+ WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14]
+ WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25]
+ WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36]
+ WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47]
+ WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58]
+ WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69]
+ WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80]
+ WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91]
+ WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101]
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110]
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119]
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] BLEQ_DN
+ BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10]
+ GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21]
+ GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32]
+ GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43]
+ GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54]
+ GW[55] GW[56] GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65]
+ GW[66] GW[67] GW[68] GW[69] GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76]
+ GW[77] GW[78] GW[79] GW[80] GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87]
+ GW[88] GW[89] GW[90] GW[91] GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98]
+ GW[99] GW[100] GW[101] GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108]
+ GW[109] GW[110] GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117]
+ GW[118] GW[119] GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126]
+ GW[127] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9]
+ GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18]
+ GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27]
+ GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36]
+ GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45]
+ GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54]
+ GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63]
+ GWB[64] GWB[65] GWB[66] GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72]
+ GWB[73] GWB[74] GWB[75] GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81]
+ GWB[82] GWB[83] GWB[84] GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90]
+ GWB[91] GWB[92] GWB[93] GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99]
+ GWB[100] GWB[101] GWB[102] GWB[103] GWB[104] GWB[105] GWB[106] GWB[107]
+ GWB[108] GWB[109] GWB[110] GWB[111] GWB[112] GWB[113] GWB[114] GWB[115]
+ GWB[116] GWB[117] GWB[118] GWB[119] GWB[120] GWB[121] GWB[122] GWB[123]
+ GWB[124] GWB[125] GWB[126] GWB[127] PREBG SAEB DEC_Y_DN[0] DEC_Y_DN[1]
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7]
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5]
+ DEC_Y_UP[6] DEC_Y_UP[7] VDDI VSSI SDBM200W80_LIO_MCB_F
XLCTRL_M_M4 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0]
+ DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6]
+ DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4]
+ DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] PREBG SAEB VDDI VSSI WLPY_DN[0] WLPY_DN[1]
+ WLPY_UP[0] WLPY_UP[1] WLP_SAE WLP_SAE_TK SDBM200W80_LCTRL_M_M4
XXDRV_STRAPD0 VDDI VSSI WLPY_DN[0] WLPY_DNB[0] SDBM200W80_XDRV_STRAP_LCNT
XXDRV_LA512_SHA_0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD0 VDDI VSSI WL[0] WL[1] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_1 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD0 VDDI VSSI WL[2] WL[3] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS1 DEC_X1[0] SH_NPD0 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_2 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD1 VDDI VSSI WL[4] WL[5] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_3 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD1 VDDI VSSI WL[6] WL[7] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS3 DEC_X1[0] SH_NPD1 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_4 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD2 VDDI VSSI WL[8] WL[9] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_5 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD2 VDDI VSSI WL[10] WL[11] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS5 DEC_X1[1] SH_NPD2 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_6 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD3 VDDI VSSI WL[12] WL[13] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_7 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD3 VDDI VSSI WL[14] WL[15] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS7 DEC_X1[1] SH_NPD3 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_8 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD4 VDDI VSSI WL[16] WL[17] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_9 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD4 VDDI VSSI WL[18] WL[19] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS9 DEC_X1[2] SH_NPD4 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_10 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD5 VDDI VSSI WL[20] WL[21] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_11 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD5 VDDI VSSI WL[22] WL[23] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS11 DEC_X1[2] SH_NPD5 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_12 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD6 VDDI VSSI WL[24] WL[25] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_13 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD6 VDDI VSSI WL[26] WL[27] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS13 DEC_X1[3] SH_NPD6 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_14 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD7 VDDI VSSI WL[28] WL[29] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_15 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD7 VDDI VSSI WL[30] WL[31] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS15 DEC_X1[3] SH_NPD7 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD8 VDDI VSSI WL[32] WL[33] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_17 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD8 VDDI VSSI WL[34] WL[35] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS17 DEC_X1[4] SH_NPD8 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_18 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD9 VDDI VSSI WL[36] WL[37] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_19 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD9 VDDI VSSI WL[38] WL[39] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS19 DEC_X1[4] SH_NPD9 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_20 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD10 VDDI VSSI WL[40] WL[41] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_21 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD10 VDDI VSSI WL[42] WL[43] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS21 DEC_X1[5] SH_NPD10 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_22 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD11 VDDI VSSI WL[44] WL[45] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_23 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD11 VDDI VSSI WL[46] WL[47] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS23 DEC_X1[5] SH_NPD11 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_24 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD12 VDDI VSSI WL[48] WL[49] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_25 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD12 VDDI VSSI WL[50] WL[51] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS25 DEC_X1[6] SH_NPD12 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_26 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD13 VDDI VSSI WL[52] WL[53] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_27 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD13 VDDI VSSI WL[54] WL[55] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS27 DEC_X1[6] SH_NPD13 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD14 VDDI VSSI WL[56] WL[57] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_29 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD14 VDDI VSSI WL[58] WL[59] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS29 DEC_X1[7] SH_NPD14 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_30 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD15 VDDI VSSI WL[60] WL[61] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_31 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD15 VDDI VSSI WL[62] WL[63] WLPY_DN[0] WLPY_DNB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS31 DEC_X1[7] SH_NPD15 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_STRAPU0 VDDI VSSI WLPY_UP[0] WLPY_UPB[0] SDBM200W80_XDRV_STRAP_LCNT
XXDRV_LA512_SHA_32 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD16 VDDI VSSI WL[64] WL[65] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_33 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD16 VDDI VSSI WL[66] WL[67] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS33 DEC_X1[0] SH_NPD16 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_34 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD17 VDDI VSSI WL[68] WL[69] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_35 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD17 VDDI VSSI WL[70] WL[71] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS35 DEC_X1[0] SH_NPD17 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_36 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD18 VDDI VSSI WL[72] WL[73] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_37 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD18 VDDI VSSI WL[74] WL[75] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS37 DEC_X1[1] SH_NPD18 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_38 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD19 VDDI VSSI WL[76] WL[77] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_39 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD19 VDDI VSSI WL[78] WL[79] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS39 DEC_X1[1] SH_NPD19 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_40 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD20 VDDI VSSI WL[80] WL[81] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_41 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD20 VDDI VSSI WL[82] WL[83] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS41 DEC_X1[2] SH_NPD20 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_42 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD21 VDDI VSSI WL[84] WL[85] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_43 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD21 VDDI VSSI WL[86] WL[87] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS43 DEC_X1[2] SH_NPD21 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_44 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD22 VDDI VSSI WL[88] WL[89] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_45 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD22 VDDI VSSI WL[90] WL[91] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS45 DEC_X1[3] SH_NPD22 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_46 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD23 VDDI VSSI WL[92] WL[93] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_47 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD23 VDDI VSSI WL[94] WL[95] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS47 DEC_X1[3] SH_NPD23 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_48 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD24 VDDI VSSI WL[96] WL[97] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_49 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD24 VDDI VSSI WL[98] WL[99] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS49 DEC_X1[4] SH_NPD24 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_50 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD25 VDDI VSSI WL[100] WL[101] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_51 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD25 VDDI VSSI WL[102] WL[103] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS51 DEC_X1[4] SH_NPD25 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_52 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD26 VDDI VSSI WL[104] WL[105] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_53 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD26 VDDI VSSI WL[106] WL[107] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS53 DEC_X1[5] SH_NPD26 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_54 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD27 VDDI VSSI WL[108] WL[109] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_55 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD27 VDDI VSSI WL[110] WL[111] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS55 DEC_X1[5] SH_NPD27 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_56 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD28 VDDI VSSI WL[112] WL[113] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_57 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD28 VDDI VSSI WL[114] WL[115] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS57 DEC_X1[6] SH_NPD28 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_58 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD29 VDDI VSSI WL[116] WL[117] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_59 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD29 VDDI VSSI WL[118] WL[119] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS59 DEC_X1[6] SH_NPD29 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_60 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD30 VDDI VSSI WL[120] WL[121] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_61 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD30 VDDI VSSI WL[122] WL[123] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS61 DEC_X1[7] SH_NPD30 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_62 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD31 VDDI VSSI WL[124] WL[125] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_63 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] SH_NPD31 VDDI VSSI WL[126] WL[127] WLPY_UP[0] WLPY_UPB[0] WLP_SAE
+ WLP_SAE_TK SDBM200W80_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS63 DEC_X1[7] SH_NPD31 VSSI SDBM200W80_XDRV_LA512_SHA_NMOS
.ENDS

.SUBCKT SDBM200W80_CNT_CORE_IO AWT AWT2 BLTRKWLDRV CEBA CEBB CKD CLK DCLKA
+ DCLK_L DCLK_R DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] DEC_X3[1]
+ DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1]
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PHASESEL_L PHASESEL_R
+ PTSEL[0] PTSEL[1] QLATCH_AB_L QLATCH_AB_R QLATCH_BB_L QLATCH_BB_R RSC_TRK_W
+ RTSEL[0] RTSEL[1] TMA TMB TRKBL VDDI VHI VLO VSSI WEBA WEBB WLP_SAE WLP_SAEB
+ WLP_SAE_TK WTSEL[0] WTSEL[1] XA[0] XA[1] XA[2] XA[3] XA[4] XA[5] XA[6] XA[7]
+ XA[8] XA[9] XB[0] XB[1] XB[2] XB[3] XB[4] XB[5] XB[6] XB[7] XB[8] XB[9] YA[0]
+ YA[1] YB[0] YB[1] BWEBA[0] BWEBA[1] BWEBA[2] BWEBA[3] BWEBA[4] BWEBA[5]
+ BWEBA[6] BWEBA[7] BWEBA[8] BWEBA[9] BWEBB[0] BWEBB[1] BWEBB[2] BWEBB[3]
+ BWEBB[4] BWEBB[5] BWEBB[6] BWEBB[7] BWEBB[8] BWEBB[9] DA[0] DA[1] DA[2] DA[3]
+ DA[4] DA[5] DA[6] DA[7] DA[8] DA[9] DB[0] DB[1] DB[2] DB[3] DB[4] DB[5] DB[6]
+ DB[7] DB[8] DB[9] GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7]
+ GBL[8] GBL[9] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7]
+ GBLB[8] GBLB[9] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] QA[0]
+ QA[1] QA[2] QA[3] QA[4] QA[5] QA[6] QA[7] QA[8] QA[9] QB[0] QB[1] QB[2] QB[3]
+ QB[4] QB[5] QB[6] QB[7] QB[8] QB[9]
XCNT_WOBIST_M4_DP_IOX10 AWT AWT2 BLTRKWLDRV BWEBA[0] BWEBA[1] BWEBA[2] BWEBA[3]
+ BWEBA[6] BWEBA[7] BWEBA[8] BWEBA[9] BWEBA[4] BWEBA[5] BWEBB[0] BWEBB[1]
+ BWEBB[2] BWEBB[3] BWEBB[6] BWEBB[7] BWEBB[8] BWEBB[9] BWEBB[4] BWEBB[5] CEBA
+ CEBB CKD CLK DA[0] DA[1] DA[2] DA[3] DA[6] DA[7] DA[8] DA[9] DA[4] DA[5] DB[0]
+ DB[1] DB[2] DB[3] DB[6] DB[7] DB[8] DB[9] DB[4] DB[5] DCLKA DCLK_L DCLK_R
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] DEC_X3[1] DEC_X3[2]
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2]
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[6] GBLB[7]
+ GBLB[8] GBLB[9] GBLB[4] GBLB[5] GBL[4] GBL[5] GW[0] GW[1] GW[2] GW[3] GW[6]
+ GW[7] GW[8] GW[9] GWB[0] GWB[1] GWB[2] GWB[3] GWB[6] GWB[7] GWB[8] GWB[9]
+ GWB[4] GWB[5] GW[4] GW[5] PHASESEL_L PHASESEL_R PTSEL[0] PTSEL[1] QA[0] QA[1]
+ QA[2] QA[3] QA[6] QA[7] QA[8] QA[9] QA[4] QA[5] QB[0] QB[1] QB[2] QB[3] QB[6]
+ QB[7] QB[8] QB[9] QB[4] QB[5] QLATCH_AB_L QLATCH_AB_R QLATCH_BB_L QLATCH_BB_R
+ RSC_TRK_W RSC_TRK_H RTSEL[0] RTSEL[1] TMA TMB TRKBL VDDI VHI VLO VSSI WEBA
+ WEBB WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] XA[0] XA[1] XA[2] XA[3]
+ XA[4] XA[5] XA[6] XA[7] XA[8] XA[9] XB[0] XB[1] XB[2] XB[3] XB[4] XB[5] XB[6]
+ XB[7] XB[8] XB[9] YA[0] YA[1] YB[0] YB[1]
+ SDBM200W80_CNT_WOBIST_M4_DP_IOX10_HALF
.ENDS

.SUBCKT SDBM200W80_MIO_L AWT BWEBA[58] BWEBA[57] BWEBA[56] BWEBA[55] BWEBA[54]
+ BWEBA[53] BWEBA[52] BWEBA[51] BWEBA[50] BWEBA[49] BWEBA[48] BWEBA[47]
+ BWEBA[46] BWEBA[45] BWEBA[44] BWEBA[43] BWEBA[42] BWEBA[41] BWEBA[40]
+ BWEBA[39] BWEBA[38] BWEBA[37] BWEBA[36] BWEBA[35] BWEBA[34] BWEBA[33]
+ BWEBA[32] BWEBA[31] BWEBA[30] BWEBA[29] BWEBA[28] BWEBA[27] BWEBA[26]
+ BWEBA[25] BWEBA[24] BWEBA[23] BWEBA[22] BWEBA[21] BWEBA[20] BWEBA[19]
+ BWEBA[18] BWEBA[17] BWEBA[16] BWEBA[15] BWEBA[14] BWEBA[13] BWEBA[12]
+ BWEBA[11] BWEBA[10] BWEBA[9] BWEBA[8] BWEBA[7] BWEBA[6] BWEBA[5] BWEBA[4]
+ BWEBA[3] BWEBA[2] BWEBA[1] BWEBA[0] BWEBB[58] BWEBB[57] BWEBB[56] BWEBB[55]
+ BWEBB[54] BWEBB[53] BWEBB[52] BWEBB[51] BWEBB[50] BWEBB[49] BWEBB[48]
+ BWEBB[47] BWEBB[46] BWEBB[45] BWEBB[44] BWEBB[43] BWEBB[42] BWEBB[41]
+ BWEBB[40] BWEBB[39] BWEBB[38] BWEBB[37] BWEBB[36] BWEBB[35] BWEBB[34]
+ BWEBB[33] BWEBB[32] BWEBB[31] BWEBB[30] BWEBB[29] BWEBB[28] BWEBB[27]
+ BWEBB[26] BWEBB[25] BWEBB[24] BWEBB[23] BWEBB[22] BWEBB[21] BWEBB[20]
+ BWEBB[19] BWEBB[18] BWEBB[17] BWEBB[16] BWEBB[15] BWEBB[14] BWEBB[13]
+ BWEBB[12] BWEBB[11] BWEBB[10] BWEBB[9] BWEBB[8] BWEBB[7] BWEBB[6] BWEBB[5]
+ BWEBB[4] BWEBB[3] BWEBB[2] BWEBB[1] BWEBB[0] CKD DA[58] DA[57] DA[56] DA[55]
+ DA[54] DA[53] DA[52] DA[51] DA[50] DA[49] DA[48] DA[47] DA[46] DA[45] DA[44]
+ DA[43] DA[42] DA[41] DA[40] DA[39] DA[38] DA[37] DA[36] DA[35] DA[34] DA[33]
+ DA[32] DA[31] DA[30] DA[29] DA[28] DA[27] DA[26] DA[25] DA[24] DA[23] DA[22]
+ DA[21] DA[20] DA[19] DA[18] DA[17] DA[16] DA[15] DA[14] DA[13] DA[12] DA[11]
+ DA[10] DA[9] DA[8] DA[7] DA[6] DA[5] DA[4] DA[3] DA[2] DA[1] DA[0] DB[58]
+ DB[57] DB[56] DB[55] DB[54] DB[53] DB[52] DB[51] DB[50] DB[49] DB[48] DB[47]
+ DB[46] DB[45] DB[44] DB[43] DB[42] DB[41] DB[40] DB[39] DB[38] DB[37] DB[36]
+ DB[35] DB[34] DB[33] DB[32] DB[31] DB[30] DB[29] DB[28] DB[27] DB[26] DB[25]
+ DB[24] DB[23] DB[22] DB[21] DB[20] DB[19] DB[18] DB[17] DB[16] DB[15] DB[14]
+ DB[13] DB[12] DB[11] DB[10] DB[9] DB[8] DB[7] DB[6] DB[5] DB[4] DB[3] DB[2]
+ DB[1] DB[0] DCLK_L DCLKA GBL[58] GBL[57] GBL[56] GBL[55] GBL[54] GBL[53]
+ GBL[52] GBL[51] GBL[50] GBL[49] GBL[48] GBL[47] GBL[46] GBL[45] GBL[44]
+ GBL[43] GBL[42] GBL[41] GBL[40] GBL[39] GBL[38] GBL[37] GBL[36] GBL[35]
+ GBL[34] GBL[33] GBL[32] GBL[31] GBL[30] GBL[29] GBL[28] GBL[27] GBL[26]
+ GBL[25] GBL[24] GBL[23] GBL[22] GBL[21] GBL[20] GBL[19] GBL[18] GBL[17]
+ GBL[16] GBL[15] GBL[14] GBL[13] GBL[12] GBL[11] GBL[10] GBL[9] GBL[8] GBL[7]
+ GBL[6] GBL[5] GBL[4] GBL[3] GBL[2] GBL[1] GBL[0] GBLB[58] GBLB[57] GBLB[56]
+ GBLB[55] GBLB[54] GBLB[53] GBLB[52] GBLB[51] GBLB[50] GBLB[49] GBLB[48]
+ GBLB[47] GBLB[46] GBLB[45] GBLB[44] GBLB[43] GBLB[42] GBLB[41] GBLB[40]
+ GBLB[39] GBLB[38] GBLB[37] GBLB[36] GBLB[35] GBLB[34] GBLB[33] GBLB[32]
+ GBLB[31] GBLB[30] GBLB[29] GBLB[28] GBLB[27] GBLB[26] GBLB[25] GBLB[24]
+ GBLB[23] GBLB[22] GBLB[21] GBLB[20] GBLB[19] GBLB[18] GBLB[17] GBLB[16]
+ GBLB[15] GBLB[14] GBLB[13] GBLB[12] GBLB[11] GBLB[10] GBLB[9] GBLB[8] GBLB[7]
+ GBLB[6] GBLB[5] GBLB[4] GBLB[3] GBLB[2] GBLB[1] GBLB[0] GW[58] GW[57] GW[56]
+ GW[55] GW[54] GW[53] GW[52] GW[51] GW[50] GW[49] GW[48] GW[47] GW[46] GW[45]
+ GW[44] GW[43] GW[42] GW[41] GW[40] GW[39] GW[38] GW[37] GW[36] GW[35] GW[34]
+ GW[33] GW[32] GW[31] GW[30] GW[29] GW[28] GW[27] GW[26] GW[25] GW[24] GW[23]
+ GW[22] GW[21] GW[20] GW[19] GW[18] GW[17] GW[16] GW[15] GW[14] GW[13] GW[12]
+ GW[11] GW[10] GW[9] GW[8] GW[7] GW[6] GW[5] GW[4] GW[3] GW[2] GW[1] GW[0]
+ GWB[58] GWB[57] GWB[56] GWB[55] GWB[54] GWB[53] GWB[52] GWB[51] GWB[50]
+ GWB[49] GWB[48] GWB[47] GWB[46] GWB[45] GWB[44] GWB[43] GWB[42] GWB[41]
+ GWB[40] GWB[39] GWB[38] GWB[37] GWB[36] GWB[35] GWB[34] GWB[33] GWB[32]
+ GWB[31] GWB[30] GWB[29] GWB[28] GWB[27] GWB[26] GWB[25] GWB[24] GWB[23]
+ GWB[22] GWB[21] GWB[20] GWB[19] GWB[18] GWB[17] GWB[16] GWB[15] GWB[14]
+ GWB[13] GWB[12] GWB[11] GWB[10] GWB[9] GWB[8] GWB[7] GWB[6] GWB[5] GWB[4]
+ GWB[3] GWB[2] GWB[1] GWB[0] PHASESEL QA[58] QA[57] QA[56] QA[55] QA[54] QA[53]
+ QA[52] QA[51] QA[50] QA[49] QA[48] QA[47] QA[46] QA[45] QA[44] QA[43] QA[42]
+ QA[41] QA[40] QA[39] QA[38] QA[37] QA[36] QA[35] QA[34] QA[33] QA[32] QA[31]
+ QA[30] QA[29] QA[28] QA[27] QA[26] QA[25] QA[24] QA[23] QA[22] QA[21] QA[20]
+ QA[19] QA[18] QA[17] QA[16] QA[15] QA[14] QA[13] QA[12] QA[11] QA[10] QA[9]
+ QA[8] QA[7] QA[6] QA[5] QA[4] QA[3] QA[2] QA[1] QA[0] QB[58] QB[57] QB[56]
+ QB[55] QB[54] QB[53] QB[52] QB[51] QB[50] QB[49] QB[48] QB[47] QB[46] QB[45]
+ QB[44] QB[43] QB[42] QB[41] QB[40] QB[39] QB[38] QB[37] QB[36] QB[35] QB[34]
+ QB[33] QB[32] QB[31] QB[30] QB[29] QB[28] QB[27] QB[26] QB[25] QB[24] QB[23]
+ QB[22] QB[21] QB[20] QB[19] QB[18] QB[17] QB[16] QB[15] QB[14] QB[13] QB[12]
+ QB[11] QB[10] QB[9] QB[8] QB[7] QB[6] QB[5] QB[4] QB[3] QB[2] QB[1] QB[0]
+ QLATCH_AB_L QLATCH_BB_L VDDI VSSI VLO WLP_SAEB
XIO_WOBIST_0 AWT BWEBA[0] BWEBB[0] CKD DA[0] DB[0] DCLK_L DCLKA GBL[0] GBLB[0]
+ GW[0] GWB[0] PHASESEL QA[0] QB[0] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_1 AWT BWEBA[1] BWEBB[1] CKD DA[1] DB[1] DCLK_L DCLKA GBL[1] GBLB[1]
+ GW[1] GWB[1] PHASESEL QA[1] QB[1] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_2 AWT BWEBA[2] BWEBB[2] CKD DA[2] DB[2] DCLK_L DCLKA GBL[2] GBLB[2]
+ GW[2] GWB[2] PHASESEL QA[2] QB[2] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_3 AWT BWEBA[3] BWEBB[3] CKD DA[3] DB[3] DCLK_L DCLKA GBL[3] GBLB[3]
+ GW[3] GWB[3] PHASESEL QA[3] QB[3] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_4 AWT BWEBA[4] BWEBB[4] CKD DA[4] DB[4] DCLK_L DCLKA GBL[4] GBLB[4]
+ GW[4] GWB[4] PHASESEL QA[4] QB[4] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_5 AWT BWEBA[5] BWEBB[5] CKD DA[5] DB[5] DCLK_L DCLKA GBL[5] GBLB[5]
+ GW[5] GWB[5] PHASESEL QA[5] QB[5] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_6 AWT BWEBA[6] BWEBB[6] CKD DA[6] DB[6] DCLK_L DCLKA GBL[6] GBLB[6]
+ GW[6] GWB[6] PHASESEL QA[6] QB[6] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_7 AWT BWEBA[7] BWEBB[7] CKD DA[7] DB[7] DCLK_L DCLKA GBL[7] GBLB[7]
+ GW[7] GWB[7] PHASESEL QA[7] QB[7] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_8 AWT BWEBA[8] BWEBB[8] CKD DA[8] DB[8] DCLK_L DCLKA GBL[8] GBLB[8]
+ GW[8] GWB[8] PHASESEL QA[8] QB[8] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_9 AWT BWEBA[9] BWEBB[9] CKD DA[9] DB[9] DCLK_L DCLKA GBL[9] GBLB[9]
+ GW[9] GWB[9] PHASESEL QA[9] QB[9] QLATCH_AB_L QLATCH_BB_L RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_10 AWT BWEBA[10] BWEBB[10] CKD DA[10] DB[10] DCLK_L DCLKA GBL[10]
+ GBLB[10] GW[10] GWB[10] PHASESEL QA[10] QB[10] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_11 AWT BWEBA[11] BWEBB[11] CKD DA[11] DB[11] DCLK_L DCLKA GBL[11]
+ GBLB[11] GW[11] GWB[11] PHASESEL QA[11] QB[11] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_12 AWT BWEBA[12] BWEBB[12] CKD DA[12] DB[12] DCLK_L DCLKA GBL[12]
+ GBLB[12] GW[12] GWB[12] PHASESEL QA[12] QB[12] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_13 AWT BWEBA[13] BWEBB[13] CKD DA[13] DB[13] DCLK_L DCLKA GBL[13]
+ GBLB[13] GW[13] GWB[13] PHASESEL QA[13] QB[13] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_14 AWT BWEBA[14] BWEBB[14] CKD DA[14] DB[14] DCLK_L DCLKA GBL[14]
+ GBLB[14] GW[14] GWB[14] PHASESEL QA[14] QB[14] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_15 AWT BWEBA[15] BWEBB[15] CKD DA[15] DB[15] DCLK_L DCLKA GBL[15]
+ GBLB[15] GW[15] GWB[15] PHASESEL QA[15] QB[15] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_16 AWT BWEBA[16] BWEBB[16] CKD DA[16] DB[16] DCLK_L DCLKA GBL[16]
+ GBLB[16] GW[16] GWB[16] PHASESEL QA[16] QB[16] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_17 AWT BWEBA[17] BWEBB[17] CKD DA[17] DB[17] DCLK_L DCLKA GBL[17]
+ GBLB[17] GW[17] GWB[17] PHASESEL QA[17] QB[17] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_18 AWT BWEBA[18] BWEBB[18] CKD DA[18] DB[18] DCLK_L DCLKA GBL[18]
+ GBLB[18] GW[18] GWB[18] PHASESEL QA[18] QB[18] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_19 AWT BWEBA[19] BWEBB[19] CKD DA[19] DB[19] DCLK_L DCLKA GBL[19]
+ GBLB[19] GW[19] GWB[19] PHASESEL QA[19] QB[19] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_20 AWT BWEBA[20] BWEBB[20] CKD DA[20] DB[20] DCLK_L DCLKA GBL[20]
+ GBLB[20] GW[20] GWB[20] PHASESEL QA[20] QB[20] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_21 AWT BWEBA[21] BWEBB[21] CKD DA[21] DB[21] DCLK_L DCLKA GBL[21]
+ GBLB[21] GW[21] GWB[21] PHASESEL QA[21] QB[21] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_22 AWT BWEBA[22] BWEBB[22] CKD DA[22] DB[22] DCLK_L DCLKA GBL[22]
+ GBLB[22] GW[22] GWB[22] PHASESEL QA[22] QB[22] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_23 AWT BWEBA[23] BWEBB[23] CKD DA[23] DB[23] DCLK_L DCLKA GBL[23]
+ GBLB[23] GW[23] GWB[23] PHASESEL QA[23] QB[23] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_24 AWT BWEBA[24] BWEBB[24] CKD DA[24] DB[24] DCLK_L DCLKA GBL[24]
+ GBLB[24] GW[24] GWB[24] PHASESEL QA[24] QB[24] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_25 AWT BWEBA[25] BWEBB[25] CKD DA[25] DB[25] DCLK_L DCLKA GBL[25]
+ GBLB[25] GW[25] GWB[25] PHASESEL QA[25] QB[25] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_26 AWT BWEBA[26] BWEBB[26] CKD DA[26] DB[26] DCLK_L DCLKA GBL[26]
+ GBLB[26] GW[26] GWB[26] PHASESEL QA[26] QB[26] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_27 AWT BWEBA[27] BWEBB[27] CKD DA[27] DB[27] DCLK_L DCLKA GBL[27]
+ GBLB[27] GW[27] GWB[27] PHASESEL QA[27] QB[27] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_28 AWT BWEBA[28] BWEBB[28] CKD DA[28] DB[28] DCLK_L DCLKA GBL[28]
+ GBLB[28] GW[28] GWB[28] PHASESEL QA[28] QB[28] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_29 AWT BWEBA[29] BWEBB[29] CKD DA[29] DB[29] DCLK_L DCLKA GBL[29]
+ GBLB[29] GW[29] GWB[29] PHASESEL QA[29] QB[29] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_30 AWT BWEBA[30] BWEBB[30] CKD DA[30] DB[30] DCLK_L DCLKA GBL[30]
+ GBLB[30] GW[30] GWB[30] PHASESEL QA[30] QB[30] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_31 AWT BWEBA[31] BWEBB[31] CKD DA[31] DB[31] DCLK_L DCLKA GBL[31]
+ GBLB[31] GW[31] GWB[31] PHASESEL QA[31] QB[31] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_32 AWT BWEBA[32] BWEBB[32] CKD DA[32] DB[32] DCLK_L DCLKA GBL[32]
+ GBLB[32] GW[32] GWB[32] PHASESEL QA[32] QB[32] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_33 AWT BWEBA[33] BWEBB[33] CKD DA[33] DB[33] DCLK_L DCLKA GBL[33]
+ GBLB[33] GW[33] GWB[33] PHASESEL QA[33] QB[33] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_34 AWT BWEBA[34] BWEBB[34] CKD DA[34] DB[34] DCLK_L DCLKA GBL[34]
+ GBLB[34] GW[34] GWB[34] PHASESEL QA[34] QB[34] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_35 AWT BWEBA[35] BWEBB[35] CKD DA[35] DB[35] DCLK_L DCLKA GBL[35]
+ GBLB[35] GW[35] GWB[35] PHASESEL QA[35] QB[35] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_36 AWT BWEBA[36] BWEBB[36] CKD DA[36] DB[36] DCLK_L DCLKA GBL[36]
+ GBLB[36] GW[36] GWB[36] PHASESEL QA[36] QB[36] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_37 AWT BWEBA[37] BWEBB[37] CKD DA[37] DB[37] DCLK_L DCLKA GBL[37]
+ GBLB[37] GW[37] GWB[37] PHASESEL QA[37] QB[37] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_38 AWT BWEBA[38] BWEBB[38] CKD DA[38] DB[38] DCLK_L DCLKA GBL[38]
+ GBLB[38] GW[38] GWB[38] PHASESEL QA[38] QB[38] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_39 AWT BWEBA[39] BWEBB[39] CKD DA[39] DB[39] DCLK_L DCLKA GBL[39]
+ GBLB[39] GW[39] GWB[39] PHASESEL QA[39] QB[39] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_40 AWT BWEBA[40] BWEBB[40] CKD DA[40] DB[40] DCLK_L DCLKA GBL[40]
+ GBLB[40] GW[40] GWB[40] PHASESEL QA[40] QB[40] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_41 AWT BWEBA[41] BWEBB[41] CKD DA[41] DB[41] DCLK_L DCLKA GBL[41]
+ GBLB[41] GW[41] GWB[41] PHASESEL QA[41] QB[41] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_42 AWT BWEBA[42] BWEBB[42] CKD DA[42] DB[42] DCLK_L DCLKA GBL[42]
+ GBLB[42] GW[42] GWB[42] PHASESEL QA[42] QB[42] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_43 AWT BWEBA[43] BWEBB[43] CKD DA[43] DB[43] DCLK_L DCLKA GBL[43]
+ GBLB[43] GW[43] GWB[43] PHASESEL QA[43] QB[43] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_44 AWT BWEBA[44] BWEBB[44] CKD DA[44] DB[44] DCLK_L DCLKA GBL[44]
+ GBLB[44] GW[44] GWB[44] PHASESEL QA[44] QB[44] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_45 AWT BWEBA[45] BWEBB[45] CKD DA[45] DB[45] DCLK_L DCLKA GBL[45]
+ GBLB[45] GW[45] GWB[45] PHASESEL QA[45] QB[45] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_46 AWT BWEBA[46] BWEBB[46] CKD DA[46] DB[46] DCLK_L DCLKA GBL[46]
+ GBLB[46] GW[46] GWB[46] PHASESEL QA[46] QB[46] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_47 AWT BWEBA[47] BWEBB[47] CKD DA[47] DB[47] DCLK_L DCLKA GBL[47]
+ GBLB[47] GW[47] GWB[47] PHASESEL QA[47] QB[47] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_48 AWT BWEBA[48] BWEBB[48] CKD DA[48] DB[48] DCLK_L DCLKA GBL[48]
+ GBLB[48] GW[48] GWB[48] PHASESEL QA[48] QB[48] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_49 AWT BWEBA[49] BWEBB[49] CKD DA[49] DB[49] DCLK_L DCLKA GBL[49]
+ GBLB[49] GW[49] GWB[49] PHASESEL QA[49] QB[49] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_50 AWT BWEBA[50] BWEBB[50] CKD DA[50] DB[50] DCLK_L DCLKA GBL[50]
+ GBLB[50] GW[50] GWB[50] PHASESEL QA[50] QB[50] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_51 AWT BWEBA[51] BWEBB[51] CKD DA[51] DB[51] DCLK_L DCLKA GBL[51]
+ GBLB[51] GW[51] GWB[51] PHASESEL QA[51] QB[51] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_52 AWT BWEBA[52] BWEBB[52] CKD DA[52] DB[52] DCLK_L DCLKA GBL[52]
+ GBLB[52] GW[52] GWB[52] PHASESEL QA[52] QB[52] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_53 AWT BWEBA[53] BWEBB[53] CKD DA[53] DB[53] DCLK_L DCLKA GBL[53]
+ GBLB[53] GW[53] GWB[53] PHASESEL QA[53] QB[53] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_54 AWT BWEBA[54] BWEBB[54] CKD DA[54] DB[54] DCLK_L DCLKA GBL[54]
+ GBLB[54] GW[54] GWB[54] PHASESEL QA[54] QB[54] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_55 AWT BWEBA[55] BWEBB[55] CKD DA[55] DB[55] DCLK_L DCLKA GBL[55]
+ GBLB[55] GW[55] GWB[55] PHASESEL QA[55] QB[55] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_56 AWT BWEBA[56] BWEBB[56] CKD DA[56] DB[56] DCLK_L DCLKA GBL[56]
+ GBLB[56] GW[56] GWB[56] PHASESEL QA[56] QB[56] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_57 AWT BWEBA[57] BWEBB[57] CKD DA[57] DB[57] DCLK_L DCLKA GBL[57]
+ GBLB[57] GW[57] GWB[57] PHASESEL QA[57] QB[57] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_58 AWT BWEBA[58] BWEBB[58] CKD DA[58] DB[58] DCLK_L DCLKA GBL[58]
+ GBLB[58] GW[58] GWB[58] PHASESEL QA[58] QB[58] QLATCH_AB_L QLATCH_BB_L
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
.ENDS

.SUBCKT SDBM200W80_MIO_R AWT BWEBA[58] BWEBA[57] BWEBA[56] BWEBA[55] BWEBA[54]
+ BWEBA[53] BWEBA[52] BWEBA[51] BWEBA[50] BWEBA[49] BWEBA[48] BWEBA[47]
+ BWEBA[46] BWEBA[45] BWEBA[44] BWEBA[43] BWEBA[42] BWEBA[41] BWEBA[40]
+ BWEBA[39] BWEBA[38] BWEBA[37] BWEBA[36] BWEBA[35] BWEBA[34] BWEBA[33]
+ BWEBA[32] BWEBA[31] BWEBA[30] BWEBA[29] BWEBA[28] BWEBA[27] BWEBA[26]
+ BWEBA[25] BWEBA[24] BWEBA[23] BWEBA[22] BWEBA[21] BWEBA[20] BWEBA[19]
+ BWEBA[18] BWEBA[17] BWEBA[16] BWEBA[15] BWEBA[14] BWEBA[13] BWEBA[12]
+ BWEBA[11] BWEBA[10] BWEBA[9] BWEBA[8] BWEBA[7] BWEBA[6] BWEBA[5] BWEBA[4]
+ BWEBA[3] BWEBA[2] BWEBA[1] BWEBA[0] BWEBB[58] BWEBB[57] BWEBB[56] BWEBB[55]
+ BWEBB[54] BWEBB[53] BWEBB[52] BWEBB[51] BWEBB[50] BWEBB[49] BWEBB[48]
+ BWEBB[47] BWEBB[46] BWEBB[45] BWEBB[44] BWEBB[43] BWEBB[42] BWEBB[41]
+ BWEBB[40] BWEBB[39] BWEBB[38] BWEBB[37] BWEBB[36] BWEBB[35] BWEBB[34]
+ BWEBB[33] BWEBB[32] BWEBB[31] BWEBB[30] BWEBB[29] BWEBB[28] BWEBB[27]
+ BWEBB[26] BWEBB[25] BWEBB[24] BWEBB[23] BWEBB[22] BWEBB[21] BWEBB[20]
+ BWEBB[19] BWEBB[18] BWEBB[17] BWEBB[16] BWEBB[15] BWEBB[14] BWEBB[13]
+ BWEBB[12] BWEBB[11] BWEBB[10] BWEBB[9] BWEBB[8] BWEBB[7] BWEBB[6] BWEBB[5]
+ BWEBB[4] BWEBB[3] BWEBB[2] BWEBB[1] BWEBB[0] CKD DA[58] DA[57] DA[56] DA[55]
+ DA[54] DA[53] DA[52] DA[51] DA[50] DA[49] DA[48] DA[47] DA[46] DA[45] DA[44]
+ DA[43] DA[42] DA[41] DA[40] DA[39] DA[38] DA[37] DA[36] DA[35] DA[34] DA[33]
+ DA[32] DA[31] DA[30] DA[29] DA[28] DA[27] DA[26] DA[25] DA[24] DA[23] DA[22]
+ DA[21] DA[20] DA[19] DA[18] DA[17] DA[16] DA[15] DA[14] DA[13] DA[12] DA[11]
+ DA[10] DA[9] DA[8] DA[7] DA[6] DA[5] DA[4] DA[3] DA[2] DA[1] DA[0] DB[58]
+ DB[57] DB[56] DB[55] DB[54] DB[53] DB[52] DB[51] DB[50] DB[49] DB[48] DB[47]
+ DB[46] DB[45] DB[44] DB[43] DB[42] DB[41] DB[40] DB[39] DB[38] DB[37] DB[36]
+ DB[35] DB[34] DB[33] DB[32] DB[31] DB[30] DB[29] DB[28] DB[27] DB[26] DB[25]
+ DB[24] DB[23] DB[22] DB[21] DB[20] DB[19] DB[18] DB[17] DB[16] DB[15] DB[14]
+ DB[13] DB[12] DB[11] DB[10] DB[9] DB[8] DB[7] DB[6] DB[5] DB[4] DB[3] DB[2]
+ DB[1] DB[0] DCLK_R DCLKA GBL[58] GBL[57] GBL[56] GBL[55] GBL[54] GBL[53]
+ GBL[52] GBL[51] GBL[50] GBL[49] GBL[48] GBL[47] GBL[46] GBL[45] GBL[44]
+ GBL[43] GBL[42] GBL[41] GBL[40] GBL[39] GBL[38] GBL[37] GBL[36] GBL[35]
+ GBL[34] GBL[33] GBL[32] GBL[31] GBL[30] GBL[29] GBL[28] GBL[27] GBL[26]
+ GBL[25] GBL[24] GBL[23] GBL[22] GBL[21] GBL[20] GBL[19] GBL[18] GBL[17]
+ GBL[16] GBL[15] GBL[14] GBL[13] GBL[12] GBL[11] GBL[10] GBL[9] GBL[8] GBL[7]
+ GBL[6] GBL[5] GBL[4] GBL[3] GBL[2] GBL[1] GBL[0] GBLB[58] GBLB[57] GBLB[56]
+ GBLB[55] GBLB[54] GBLB[53] GBLB[52] GBLB[51] GBLB[50] GBLB[49] GBLB[48]
+ GBLB[47] GBLB[46] GBLB[45] GBLB[44] GBLB[43] GBLB[42] GBLB[41] GBLB[40]
+ GBLB[39] GBLB[38] GBLB[37] GBLB[36] GBLB[35] GBLB[34] GBLB[33] GBLB[32]
+ GBLB[31] GBLB[30] GBLB[29] GBLB[28] GBLB[27] GBLB[26] GBLB[25] GBLB[24]
+ GBLB[23] GBLB[22] GBLB[21] GBLB[20] GBLB[19] GBLB[18] GBLB[17] GBLB[16]
+ GBLB[15] GBLB[14] GBLB[13] GBLB[12] GBLB[11] GBLB[10] GBLB[9] GBLB[8] GBLB[7]
+ GBLB[6] GBLB[5] GBLB[4] GBLB[3] GBLB[2] GBLB[1] GBLB[0] GW[58] GW[57] GW[56]
+ GW[55] GW[54] GW[53] GW[52] GW[51] GW[50] GW[49] GW[48] GW[47] GW[46] GW[45]
+ GW[44] GW[43] GW[42] GW[41] GW[40] GW[39] GW[38] GW[37] GW[36] GW[35] GW[34]
+ GW[33] GW[32] GW[31] GW[30] GW[29] GW[28] GW[27] GW[26] GW[25] GW[24] GW[23]
+ GW[22] GW[21] GW[20] GW[19] GW[18] GW[17] GW[16] GW[15] GW[14] GW[13] GW[12]
+ GW[11] GW[10] GW[9] GW[8] GW[7] GW[6] GW[5] GW[4] GW[3] GW[2] GW[1] GW[0]
+ GWB[58] GWB[57] GWB[56] GWB[55] GWB[54] GWB[53] GWB[52] GWB[51] GWB[50]
+ GWB[49] GWB[48] GWB[47] GWB[46] GWB[45] GWB[44] GWB[43] GWB[42] GWB[41]
+ GWB[40] GWB[39] GWB[38] GWB[37] GWB[36] GWB[35] GWB[34] GWB[33] GWB[32]
+ GWB[31] GWB[30] GWB[29] GWB[28] GWB[27] GWB[26] GWB[25] GWB[24] GWB[23]
+ GWB[22] GWB[21] GWB[20] GWB[19] GWB[18] GWB[17] GWB[16] GWB[15] GWB[14]
+ GWB[13] GWB[12] GWB[11] GWB[10] GWB[9] GWB[8] GWB[7] GWB[6] GWB[5] GWB[4]
+ GWB[3] GWB[2] GWB[1] GWB[0] PHASESEL QA[58] QA[57] QA[56] QA[55] QA[54] QA[53]
+ QA[52] QA[51] QA[50] QA[49] QA[48] QA[47] QA[46] QA[45] QA[44] QA[43] QA[42]
+ QA[41] QA[40] QA[39] QA[38] QA[37] QA[36] QA[35] QA[34] QA[33] QA[32] QA[31]
+ QA[30] QA[29] QA[28] QA[27] QA[26] QA[25] QA[24] QA[23] QA[22] QA[21] QA[20]
+ QA[19] QA[18] QA[17] QA[16] QA[15] QA[14] QA[13] QA[12] QA[11] QA[10] QA[9]
+ QA[8] QA[7] QA[6] QA[5] QA[4] QA[3] QA[2] QA[1] QA[0] QB[58] QB[57] QB[56]
+ QB[55] QB[54] QB[53] QB[52] QB[51] QB[50] QB[49] QB[48] QB[47] QB[46] QB[45]
+ QB[44] QB[43] QB[42] QB[41] QB[40] QB[39] QB[38] QB[37] QB[36] QB[35] QB[34]
+ QB[33] QB[32] QB[31] QB[30] QB[29] QB[28] QB[27] QB[26] QB[25] QB[24] QB[23]
+ QB[22] QB[21] QB[20] QB[19] QB[18] QB[17] QB[16] QB[15] QB[14] QB[13] QB[12]
+ QB[11] QB[10] QB[9] QB[8] QB[7] QB[6] QB[5] QB[4] QB[3] QB[2] QB[1] QB[0]
+ QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI VLO WLP_SAEB
XIO_WOBIST_0 AWT BWEBA[0] BWEBB[0] CKD DA[0] DB[0] DCLK_R DCLKA GBL[0] GBLB[0]
+ GW[0] GWB[0] PHASESEL QA[0] QB[0] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_1 AWT BWEBA[1] BWEBB[1] CKD DA[1] DB[1] DCLK_R DCLKA GBL[1] GBLB[1]
+ GW[1] GWB[1] PHASESEL QA[1] QB[1] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_2 AWT BWEBA[2] BWEBB[2] CKD DA[2] DB[2] DCLK_R DCLKA GBL[2] GBLB[2]
+ GW[2] GWB[2] PHASESEL QA[2] QB[2] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_3 AWT BWEBA[3] BWEBB[3] CKD DA[3] DB[3] DCLK_R DCLKA GBL[3] GBLB[3]
+ GW[3] GWB[3] PHASESEL QA[3] QB[3] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_4 AWT BWEBA[4] BWEBB[4] CKD DA[4] DB[4] DCLK_R DCLKA GBL[4] GBLB[4]
+ GW[4] GWB[4] PHASESEL QA[4] QB[4] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_5 AWT BWEBA[5] BWEBB[5] CKD DA[5] DB[5] DCLK_R DCLKA GBL[5] GBLB[5]
+ GW[5] GWB[5] PHASESEL QA[5] QB[5] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_6 AWT BWEBA[6] BWEBB[6] CKD DA[6] DB[6] DCLK_R DCLKA GBL[6] GBLB[6]
+ GW[6] GWB[6] PHASESEL QA[6] QB[6] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_7 AWT BWEBA[7] BWEBB[7] CKD DA[7] DB[7] DCLK_R DCLKA GBL[7] GBLB[7]
+ GW[7] GWB[7] PHASESEL QA[7] QB[7] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_8 AWT BWEBA[8] BWEBB[8] CKD DA[8] DB[8] DCLK_R DCLKA GBL[8] GBLB[8]
+ GW[8] GWB[8] PHASESEL QA[8] QB[8] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_9 AWT BWEBA[9] BWEBB[9] CKD DA[9] DB[9] DCLK_R DCLKA GBL[9] GBLB[9]
+ GW[9] GWB[9] PHASESEL QA[9] QB[9] QLATCH_AB_R QLATCH_BB_R RSC_TRK_W VDDI VSSI
+ WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_10 AWT BWEBA[10] BWEBB[10] CKD DA[10] DB[10] DCLK_R DCLKA GBL[10]
+ GBLB[10] GW[10] GWB[10] PHASESEL QA[10] QB[10] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_11 AWT BWEBA[11] BWEBB[11] CKD DA[11] DB[11] DCLK_R DCLKA GBL[11]
+ GBLB[11] GW[11] GWB[11] PHASESEL QA[11] QB[11] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_12 AWT BWEBA[12] BWEBB[12] CKD DA[12] DB[12] DCLK_R DCLKA GBL[12]
+ GBLB[12] GW[12] GWB[12] PHASESEL QA[12] QB[12] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_13 AWT BWEBA[13] BWEBB[13] CKD DA[13] DB[13] DCLK_R DCLKA GBL[13]
+ GBLB[13] GW[13] GWB[13] PHASESEL QA[13] QB[13] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_14 AWT BWEBA[14] BWEBB[14] CKD DA[14] DB[14] DCLK_R DCLKA GBL[14]
+ GBLB[14] GW[14] GWB[14] PHASESEL QA[14] QB[14] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_15 AWT BWEBA[15] BWEBB[15] CKD DA[15] DB[15] DCLK_R DCLKA GBL[15]
+ GBLB[15] GW[15] GWB[15] PHASESEL QA[15] QB[15] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_16 AWT BWEBA[16] BWEBB[16] CKD DA[16] DB[16] DCLK_R DCLKA GBL[16]
+ GBLB[16] GW[16] GWB[16] PHASESEL QA[16] QB[16] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_17 AWT BWEBA[17] BWEBB[17] CKD DA[17] DB[17] DCLK_R DCLKA GBL[17]
+ GBLB[17] GW[17] GWB[17] PHASESEL QA[17] QB[17] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_18 AWT BWEBA[18] BWEBB[18] CKD DA[18] DB[18] DCLK_R DCLKA GBL[18]
+ GBLB[18] GW[18] GWB[18] PHASESEL QA[18] QB[18] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_19 AWT BWEBA[19] BWEBB[19] CKD DA[19] DB[19] DCLK_R DCLKA GBL[19]
+ GBLB[19] GW[19] GWB[19] PHASESEL QA[19] QB[19] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_20 AWT BWEBA[20] BWEBB[20] CKD DA[20] DB[20] DCLK_R DCLKA GBL[20]
+ GBLB[20] GW[20] GWB[20] PHASESEL QA[20] QB[20] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_21 AWT BWEBA[21] BWEBB[21] CKD DA[21] DB[21] DCLK_R DCLKA GBL[21]
+ GBLB[21] GW[21] GWB[21] PHASESEL QA[21] QB[21] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_22 AWT BWEBA[22] BWEBB[22] CKD DA[22] DB[22] DCLK_R DCLKA GBL[22]
+ GBLB[22] GW[22] GWB[22] PHASESEL QA[22] QB[22] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_23 AWT BWEBA[23] BWEBB[23] CKD DA[23] DB[23] DCLK_R DCLKA GBL[23]
+ GBLB[23] GW[23] GWB[23] PHASESEL QA[23] QB[23] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_24 AWT BWEBA[24] BWEBB[24] CKD DA[24] DB[24] DCLK_R DCLKA GBL[24]
+ GBLB[24] GW[24] GWB[24] PHASESEL QA[24] QB[24] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_25 AWT BWEBA[25] BWEBB[25] CKD DA[25] DB[25] DCLK_R DCLKA GBL[25]
+ GBLB[25] GW[25] GWB[25] PHASESEL QA[25] QB[25] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_26 AWT BWEBA[26] BWEBB[26] CKD DA[26] DB[26] DCLK_R DCLKA GBL[26]
+ GBLB[26] GW[26] GWB[26] PHASESEL QA[26] QB[26] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_27 AWT BWEBA[27] BWEBB[27] CKD DA[27] DB[27] DCLK_R DCLKA GBL[27]
+ GBLB[27] GW[27] GWB[27] PHASESEL QA[27] QB[27] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_28 AWT BWEBA[28] BWEBB[28] CKD DA[28] DB[28] DCLK_R DCLKA GBL[28]
+ GBLB[28] GW[28] GWB[28] PHASESEL QA[28] QB[28] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_29 AWT BWEBA[29] BWEBB[29] CKD DA[29] DB[29] DCLK_R DCLKA GBL[29]
+ GBLB[29] GW[29] GWB[29] PHASESEL QA[29] QB[29] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_30 AWT BWEBA[30] BWEBB[30] CKD DA[30] DB[30] DCLK_R DCLKA GBL[30]
+ GBLB[30] GW[30] GWB[30] PHASESEL QA[30] QB[30] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_31 AWT BWEBA[31] BWEBB[31] CKD DA[31] DB[31] DCLK_R DCLKA GBL[31]
+ GBLB[31] GW[31] GWB[31] PHASESEL QA[31] QB[31] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_32 AWT BWEBA[32] BWEBB[32] CKD DA[32] DB[32] DCLK_R DCLKA GBL[32]
+ GBLB[32] GW[32] GWB[32] PHASESEL QA[32] QB[32] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_33 AWT BWEBA[33] BWEBB[33] CKD DA[33] DB[33] DCLK_R DCLKA GBL[33]
+ GBLB[33] GW[33] GWB[33] PHASESEL QA[33] QB[33] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_34 AWT BWEBA[34] BWEBB[34] CKD DA[34] DB[34] DCLK_R DCLKA GBL[34]
+ GBLB[34] GW[34] GWB[34] PHASESEL QA[34] QB[34] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_35 AWT BWEBA[35] BWEBB[35] CKD DA[35] DB[35] DCLK_R DCLKA GBL[35]
+ GBLB[35] GW[35] GWB[35] PHASESEL QA[35] QB[35] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_36 AWT BWEBA[36] BWEBB[36] CKD DA[36] DB[36] DCLK_R DCLKA GBL[36]
+ GBLB[36] GW[36] GWB[36] PHASESEL QA[36] QB[36] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_37 AWT BWEBA[37] BWEBB[37] CKD DA[37] DB[37] DCLK_R DCLKA GBL[37]
+ GBLB[37] GW[37] GWB[37] PHASESEL QA[37] QB[37] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_38 AWT BWEBA[38] BWEBB[38] CKD DA[38] DB[38] DCLK_R DCLKA GBL[38]
+ GBLB[38] GW[38] GWB[38] PHASESEL QA[38] QB[38] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_39 AWT BWEBA[39] BWEBB[39] CKD DA[39] DB[39] DCLK_R DCLKA GBL[39]
+ GBLB[39] GW[39] GWB[39] PHASESEL QA[39] QB[39] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_40 AWT BWEBA[40] BWEBB[40] CKD DA[40] DB[40] DCLK_R DCLKA GBL[40]
+ GBLB[40] GW[40] GWB[40] PHASESEL QA[40] QB[40] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_41 AWT BWEBA[41] BWEBB[41] CKD DA[41] DB[41] DCLK_R DCLKA GBL[41]
+ GBLB[41] GW[41] GWB[41] PHASESEL QA[41] QB[41] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_42 AWT BWEBA[42] BWEBB[42] CKD DA[42] DB[42] DCLK_R DCLKA GBL[42]
+ GBLB[42] GW[42] GWB[42] PHASESEL QA[42] QB[42] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_43 AWT BWEBA[43] BWEBB[43] CKD DA[43] DB[43] DCLK_R DCLKA GBL[43]
+ GBLB[43] GW[43] GWB[43] PHASESEL QA[43] QB[43] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_44 AWT BWEBA[44] BWEBB[44] CKD DA[44] DB[44] DCLK_R DCLKA GBL[44]
+ GBLB[44] GW[44] GWB[44] PHASESEL QA[44] QB[44] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_45 AWT BWEBA[45] BWEBB[45] CKD DA[45] DB[45] DCLK_R DCLKA GBL[45]
+ GBLB[45] GW[45] GWB[45] PHASESEL QA[45] QB[45] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_46 AWT BWEBA[46] BWEBB[46] CKD DA[46] DB[46] DCLK_R DCLKA GBL[46]
+ GBLB[46] GW[46] GWB[46] PHASESEL QA[46] QB[46] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_47 AWT BWEBA[47] BWEBB[47] CKD DA[47] DB[47] DCLK_R DCLKA GBL[47]
+ GBLB[47] GW[47] GWB[47] PHASESEL QA[47] QB[47] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_48 AWT BWEBA[48] BWEBB[48] CKD DA[48] DB[48] DCLK_R DCLKA GBL[48]
+ GBLB[48] GW[48] GWB[48] PHASESEL QA[48] QB[48] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_49 AWT BWEBA[49] BWEBB[49] CKD DA[49] DB[49] DCLK_R DCLKA GBL[49]
+ GBLB[49] GW[49] GWB[49] PHASESEL QA[49] QB[49] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_50 AWT BWEBA[50] BWEBB[50] CKD DA[50] DB[50] DCLK_R DCLKA GBL[50]
+ GBLB[50] GW[50] GWB[50] PHASESEL QA[50] QB[50] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_51 AWT BWEBA[51] BWEBB[51] CKD DA[51] DB[51] DCLK_R DCLKA GBL[51]
+ GBLB[51] GW[51] GWB[51] PHASESEL QA[51] QB[51] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_52 AWT BWEBA[52] BWEBB[52] CKD DA[52] DB[52] DCLK_R DCLKA GBL[52]
+ GBLB[52] GW[52] GWB[52] PHASESEL QA[52] QB[52] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_53 AWT BWEBA[53] BWEBB[53] CKD DA[53] DB[53] DCLK_R DCLKA GBL[53]
+ GBLB[53] GW[53] GWB[53] PHASESEL QA[53] QB[53] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_54 AWT BWEBA[54] BWEBB[54] CKD DA[54] DB[54] DCLK_R DCLKA GBL[54]
+ GBLB[54] GW[54] GWB[54] PHASESEL QA[54] QB[54] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_55 AWT BWEBA[55] BWEBB[55] CKD DA[55] DB[55] DCLK_R DCLKA GBL[55]
+ GBLB[55] GW[55] GWB[55] PHASESEL QA[55] QB[55] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_56 AWT BWEBA[56] BWEBB[56] CKD DA[56] DB[56] DCLK_R DCLKA GBL[56]
+ GBLB[56] GW[56] GWB[56] PHASESEL QA[56] QB[56] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_57 AWT BWEBA[57] BWEBB[57] CKD DA[57] DB[57] DCLK_R DCLKA GBL[57]
+ GBLB[57] GW[57] GWB[57] PHASESEL QA[57] QB[57] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
XIO_WOBIST_58 AWT BWEBA[58] BWEBB[58] CKD DA[58] DB[58] DCLK_R DCLKA GBL[58]
+ GBLB[58] GW[58] GWB[58] PHASESEL QA[58] QB[58] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDDI VSSI WLP_SAEB SDBM200W80_IO_WOBIST_DP
.ENDS

.SUBCKT TSDN28HPCPUHDB512X128M4M QA[0] QA[1] QA[2] QA[3] QA[4] QA[5] QA[6] QA[7]
+ QA[8] QA[9] QA[10] QA[11] QA[12] QA[13] QA[14] QA[15] QA[16] QA[17] QA[18]
+ QA[19] QA[20] QA[21] QA[22] QA[23] QA[24] QA[25] QA[26] QA[27] QA[28] QA[29]
+ QA[30] QA[31] QA[32] QA[33] QA[34] QA[35] QA[36] QA[37] QA[38] QA[39] QA[40]
+ QA[41] QA[42] QA[43] QA[44] QA[45] QA[46] QA[47] QA[48] QA[49] QA[50] QA[51]
+ QA[52] QA[53] QA[54] QA[55] QA[56] QA[57] QA[58] QA[59] QA[60] QA[61] QA[62]
+ QA[63] QA[64] QA[65] QA[66] QA[67] QA[68] QA[69] QA[70] QA[71] QA[72] QA[73]
+ QA[74] QA[75] QA[76] QA[77] QA[78] QA[79] QA[80] QA[81] QA[82] QA[83] QA[84]
+ QA[85] QA[86] QA[87] QA[88] QA[89] QA[90] QA[91] QA[92] QA[93] QA[94] QA[95]
+ QA[96] QA[97] QA[98] QA[99] QA[100] QA[101] QA[102] QA[103] QA[104] QA[105]
+ QA[106] QA[107] QA[108] QA[109] QA[110] QA[111] QA[112] QA[113] QA[114]
+ QA[115] QA[116] QA[117] QA[118] QA[119] QA[120] QA[121] QA[122] QA[123]
+ QA[124] QA[125] QA[126] QA[127] QB[0] QB[1] QB[2] QB[3] QB[4] QB[5] QB[6]
+ QB[7] QB[8] QB[9] QB[10] QB[11] QB[12] QB[13] QB[14] QB[15] QB[16] QB[17]
+ QB[18] QB[19] QB[20] QB[21] QB[22] QB[23] QB[24] QB[25] QB[26] QB[27] QB[28]
+ QB[29] QB[30] QB[31] QB[32] QB[33] QB[34] QB[35] QB[36] QB[37] QB[38] QB[39]
+ QB[40] QB[41] QB[42] QB[43] QB[44] QB[45] QB[46] QB[47] QB[48] QB[49] QB[50]
+ QB[51] QB[52] QB[53] QB[54] QB[55] QB[56] QB[57] QB[58] QB[59] QB[60] QB[61]
+ QB[62] QB[63] QB[64] QB[65] QB[66] QB[67] QB[68] QB[69] QB[70] QB[71] QB[72]
+ QB[73] QB[74] QB[75] QB[76] QB[77] QB[78] QB[79] QB[80] QB[81] QB[82] QB[83]
+ QB[84] QB[85] QB[86] QB[87] QB[88] QB[89] QB[90] QB[91] QB[92] QB[93] QB[94]
+ QB[95] QB[96] QB[97] QB[98] QB[99] QB[100] QB[101] QB[102] QB[103] QB[104]
+ QB[105] QB[106] QB[107] QB[108] QB[109] QB[110] QB[111] QB[112] QB[113]
+ QB[114] QB[115] QB[116] QB[117] QB[118] QB[119] QB[120] QB[121] QB[122]
+ QB[123] QB[124] QB[125] QB[126] QB[127] AA[0] AA[1] AA[2] AA[3] AA[4] AA[5]
+ AA[6] AA[7] AA[8] AB[0] AB[1] AB[2] AB[3] AB[4] AB[5] AB[6] AB[7] AB[8] CEBA
+ CEBB CLK DB[0] DB[1] DB[2] DB[3] DB[4] DB[5] DB[6] DB[7] DB[8] DB[9] DB[10]
+ DB[11] DB[12] DB[13] DB[14] DB[15] DB[16] DB[17] DB[18] DB[19] DB[20] DB[21]
+ DB[22] DB[23] DB[24] DB[25] DB[26] DB[27] DB[28] DB[29] DB[30] DB[31] DB[32]
+ DB[33] DB[34] DB[35] DB[36] DB[37] DB[38] DB[39] DB[40] DB[41] DB[42] DB[43]
+ DB[44] DB[45] DB[46] DB[47] DB[48] DB[49] DB[50] DB[51] DB[52] DB[53] DB[54]
+ DB[55] DB[56] DB[57] DB[58] DB[59] DB[60] DB[61] DB[62] DB[63] DB[64] DB[65]
+ DB[66] DB[67] DB[68] DB[69] DB[70] DB[71] DB[72] DB[73] DB[74] DB[75] DB[76]
+ DB[77] DB[78] DB[79] DB[80] DB[81] DB[82] DB[83] DB[84] DB[85] DB[86] DB[87]
+ DB[88] DB[89] DB[90] DB[91] DB[92] DB[93] DB[94] DB[95] DB[96] DB[97] DB[98]
+ DB[99] DB[100] DB[101] DB[102] DB[103] DB[104] DB[105] DB[106] DB[107] DB[108]
+ DB[109] DB[110] DB[111] DB[112] DB[113] DB[114] DB[115] DB[116] DB[117]
+ DB[118] DB[119] DB[120] DB[121] DB[122] DB[123] DB[124] DB[125] DB[126]
+ DB[127] DA[0] DA[1] DA[2] DA[3] DA[4] DA[5] DA[6] DA[7] DA[8] DA[9] DA[10]
+ DA[11] DA[12] DA[13] DA[14] DA[15] DA[16] DA[17] DA[18] DA[19] DA[20] DA[21]
+ DA[22] DA[23] DA[24] DA[25] DA[26] DA[27] DA[28] DA[29] DA[30] DA[31] DA[32]
+ DA[33] DA[34] DA[35] DA[36] DA[37] DA[38] DA[39] DA[40] DA[41] DA[42] DA[43]
+ DA[44] DA[45] DA[46] DA[47] DA[48] DA[49] DA[50] DA[51] DA[52] DA[53] DA[54]
+ DA[55] DA[56] DA[57] DA[58] DA[59] DA[60] DA[61] DA[62] DA[63] DA[64] DA[65]
+ DA[66] DA[67] DA[68] DA[69] DA[70] DA[71] DA[72] DA[73] DA[74] DA[75] DA[76]
+ DA[77] DA[78] DA[79] DA[80] DA[81] DA[82] DA[83] DA[84] DA[85] DA[86] DA[87]
+ DA[88] DA[89] DA[90] DA[91] DA[92] DA[93] DA[94] DA[95] DA[96] DA[97] DA[98]
+ DA[99] DA[100] DA[101] DA[102] DA[103] DA[104] DA[105] DA[106] DA[107] DA[108]
+ DA[109] DA[110] DA[111] DA[112] DA[113] DA[114] DA[115] DA[116] DA[117]
+ DA[118] DA[119] DA[120] DA[121] DA[122] DA[123] DA[124] DA[125] DA[126]
+ DA[127] RTSEL[0] RTSEL[1] PTSEL[0] PTSEL[1] WTSEL[0] WTSEL[1] WEBA WEBB VDD
+ VSS
XBANK_0 GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36]
+ GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45]
+ GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54]
+ GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63]
+ GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBL[69] GBL[70] GBL[71] GBL[72]
+ GBL[73] GBL[74] GBL[75] GBL[76] GBL[77] GBL[78] GBL[79] GBL[80] GBL[81]
+ GBL[82] GBL[83] GBL[84] GBL[85] GBL[86] GBL[87] GBL[88] GBL[89] GBL[90]
+ GBL[91] GBL[92] GBL[93] GBL[94] GBL[95] GBL[96] GBL[97] GBL[98] GBL[99]
+ GBL[100] GBL[101] GBL[102] GBL[103] GBL[104] GBL[105] GBL[106] GBL[107]
+ GBL[108] GBL[109] GBL[110] GBL[111] GBL[112] GBL[113] GBL[114] GBL[115]
+ GBL[116] GBL[117] GBL[118] GBL[119] GBL[120] GBL[121] GBL[122] GBL[123]
+ GBL[124] GBL[125] GBL[126] GBL[127] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37]
+ GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45]
+ GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53]
+ GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61]
+ GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67] GBLB[68] GBLB[69]
+ GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75] GBLB[76] GBLB[77]
+ GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83] GBLB[84] GBLB[85]
+ GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91] GBLB[92] GBLB[93]
+ GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99] GBLB[100] GBLB[101]
+ GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106] GBLB[107] GBLB[108]
+ GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113] GBLB[114] GBLB[115]
+ GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120] GBLB[121] GBLB[122]
+ GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67] GW[68] GW[69] GW[70]
+ GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78] GW[79] GW[80] GW[81]
+ GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89] GW[90] GW[91] GW[92]
+ GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100] GW[101] GW[102]
+ GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109] GW[110] GW[111]
+ GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118] GW[119] GW[120]
+ GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[0] GWB[1] GWB[2]
+ GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12]
+ GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21]
+ GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30]
+ GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39]
+ GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48]
+ GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57]
+ GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65] GWB[66]
+ GWB[67] GWB[68] GWB[69] GWB[70] GWB[71] GWB[72] GWB[73] GWB[74] GWB[75]
+ GWB[76] GWB[77] GWB[78] GWB[79] GWB[80] GWB[81] GWB[82] GWB[83] GWB[84]
+ GWB[85] GWB[86] GWB[87] GWB[88] GWB[89] GWB[90] GWB[91] GWB[92] GWB[93]
+ GWB[94] GWB[95] GWB[96] GWB[97] GWB[98] GWB[99] GWB[100] GWB[101] GWB[102]
+ GWB[103] GWB[104] GWB[105] GWB[106] GWB[107] GWB[108] GWB[109] GWB[110]
+ GWB[111] GWB[112] GWB[113] GWB[114] GWB[115] GWB[116] GWB[117] GWB[118]
+ GWB[119] GWB[120] GWB[121] GWB[122] GWB[123] GWB[124] GWB[125] GWB[126]
+ GWB[127] SLP_LCTRL WLP_SAE DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] TRKBL BLTRKWLDRV VDD VSS WLP_SAE_TK SDBM200W80_BANK_0_F
XMIO_L AWT2 VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO CKD DA[0] DA[1] DA[2] DA[3] DA[4] DA[5] DA[6] DA[7]
+ DA[8] DA[9] DA[10] DA[11] DA[12] DA[13] DA[14] DA[15] DA[16] DA[17] DA[18]
+ DA[19] DA[20] DA[21] DA[22] DA[23] DA[24] DA[25] DA[26] DA[27] DA[28] DA[29]
+ DA[30] DA[31] DA[32] DA[33] DA[34] DA[35] DA[36] DA[37] DA[38] DA[39] DA[40]
+ DA[41] DA[42] DA[43] DA[44] DA[45] DA[46] DA[47] DA[48] DA[49] DA[50] DA[51]
+ DA[52] DA[53] DA[54] DA[55] DA[56] DA[57] DA[58] DB[0] DB[1] DB[2] DB[3] DB[4]
+ DB[5] DB[6] DB[7] DB[8] DB[9] DB[10] DB[11] DB[12] DB[13] DB[14] DB[15] DB[16]
+ DB[17] DB[18] DB[19] DB[20] DB[21] DB[22] DB[23] DB[24] DB[25] DB[26] DB[27]
+ DB[28] DB[29] DB[30] DB[31] DB[32] DB[33] DB[34] DB[35] DB[36] DB[37] DB[38]
+ DB[39] DB[40] DB[41] DB[42] DB[43] DB[44] DB[45] DB[46] DB[47] DB[48] DB[49]
+ DB[50] DB[51] DB[52] DB[53] DB[54] DB[55] DB[56] DB[57] DB[58] DCLK_L DCLKA
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5]
+ GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14]
+ GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22]
+ GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30]
+ GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38]
+ GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46]
+ GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54]
+ GBLB[55] GBLB[56] GBLB[57] GBLB[58] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6]
+ GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17]
+ GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28]
+ GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39]
+ GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50]
+ GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GWB[0] GWB[1] GWB[2]
+ GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12]
+ GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21]
+ GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30]
+ GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39]
+ GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48]
+ GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57]
+ GWB[58] PHASESEL_L QA[0] QA[1] QA[2] QA[3] QA[4] QA[5] QA[6] QA[7] QA[8] QA[9]
+ QA[10] QA[11] QA[12] QA[13] QA[14] QA[15] QA[16] QA[17] QA[18] QA[19] QA[20]
+ QA[21] QA[22] QA[23] QA[24] QA[25] QA[26] QA[27] QA[28] QA[29] QA[30] QA[31]
+ QA[32] QA[33] QA[34] QA[35] QA[36] QA[37] QA[38] QA[39] QA[40] QA[41] QA[42]
+ QA[43] QA[44] QA[45] QA[46] QA[47] QA[48] QA[49] QA[50] QA[51] QA[52] QA[53]
+ QA[54] QA[55] QA[56] QA[57] QA[58] QB[0] QB[1] QB[2] QB[3] QB[4] QB[5] QB[6]
+ QB[7] QB[8] QB[9] QB[10] QB[11] QB[12] QB[13] QB[14] QB[15] QB[16] QB[17]
+ QB[18] QB[19] QB[20] QB[21] QB[22] QB[23] QB[24] QB[25] QB[26] QB[27] QB[28]
+ QB[29] QB[30] QB[31] QB[32] QB[33] QB[34] QB[35] QB[36] QB[37] QB[38] QB[39]
+ QB[40] QB[41] QB[42] QB[43] QB[44] QB[45] QB[46] QB[47] QB[48] QB[49] QB[50]
+ QB[51] QB[52] QB[53] QB[54] QB[55] QB[56] QB[57] QB[58] QLATCH_AB_L
+ QLATCH_BB_L VDD VSS VLO WLP_SAEB SDBM200W80_MIO_L
XMIO_R AWT2 VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ VLO VLO VLO VLO VLO VLO CKD DA[69] DA[70] DA[71] DA[72] DA[73] DA[74] DA[75]
+ DA[76] DA[77] DA[78] DA[79] DA[80] DA[81] DA[82] DA[83] DA[84] DA[85] DA[86]
+ DA[87] DA[88] DA[89] DA[90] DA[91] DA[92] DA[93] DA[94] DA[95] DA[96] DA[97]
+ DA[98] DA[99] DA[100] DA[101] DA[102] DA[103] DA[104] DA[105] DA[106] DA[107]
+ DA[108] DA[109] DA[110] DA[111] DA[112] DA[113] DA[114] DA[115] DA[116]
+ DA[117] DA[118] DA[119] DA[120] DA[121] DA[122] DA[123] DA[124] DA[125]
+ DA[126] DA[127] DB[69] DB[70] DB[71] DB[72] DB[73] DB[74] DB[75] DB[76] DB[77]
+ DB[78] DB[79] DB[80] DB[81] DB[82] DB[83] DB[84] DB[85] DB[86] DB[87] DB[88]
+ DB[89] DB[90] DB[91] DB[92] DB[93] DB[94] DB[95] DB[96] DB[97] DB[98] DB[99]
+ DB[100] DB[101] DB[102] DB[103] DB[104] DB[105] DB[106] DB[107] DB[108]
+ DB[109] DB[110] DB[111] DB[112] DB[113] DB[114] DB[115] DB[116] DB[117]
+ DB[118] DB[119] DB[120] DB[121] DB[122] DB[123] DB[124] DB[125] DB[126]
+ DB[127] DCLK_R DCLKA GBL[69] GBL[70] GBL[71] GBL[72] GBL[73] GBL[74] GBL[75]
+ GBL[76] GBL[77] GBL[78] GBL[79] GBL[80] GBL[81] GBL[82] GBL[83] GBL[84]
+ GBL[85] GBL[86] GBL[87] GBL[88] GBL[89] GBL[90] GBL[91] GBL[92] GBL[93]
+ GBL[94] GBL[95] GBL[96] GBL[97] GBL[98] GBL[99] GBL[100] GBL[101] GBL[102]
+ GBL[103] GBL[104] GBL[105] GBL[106] GBL[107] GBL[108] GBL[109] GBL[110]
+ GBL[111] GBL[112] GBL[113] GBL[114] GBL[115] GBL[116] GBL[117] GBL[118]
+ GBL[119] GBL[120] GBL[121] GBL[122] GBL[123] GBL[124] GBL[125] GBL[126]
+ GBL[127] GBLB[69] GBLB[70] GBLB[71] GBLB[72] GBLB[73] GBLB[74] GBLB[75]
+ GBLB[76] GBLB[77] GBLB[78] GBLB[79] GBLB[80] GBLB[81] GBLB[82] GBLB[83]
+ GBLB[84] GBLB[85] GBLB[86] GBLB[87] GBLB[88] GBLB[89] GBLB[90] GBLB[91]
+ GBLB[92] GBLB[93] GBLB[94] GBLB[95] GBLB[96] GBLB[97] GBLB[98] GBLB[99]
+ GBLB[100] GBLB[101] GBLB[102] GBLB[103] GBLB[104] GBLB[105] GBLB[106]
+ GBLB[107] GBLB[108] GBLB[109] GBLB[110] GBLB[111] GBLB[112] GBLB[113]
+ GBLB[114] GBLB[115] GBLB[116] GBLB[117] GBLB[118] GBLB[119] GBLB[120]
+ GBLB[121] GBLB[122] GBLB[123] GBLB[124] GBLB[125] GBLB[126] GBLB[127] GW[69]
+ GW[70] GW[71] GW[72] GW[73] GW[74] GW[75] GW[76] GW[77] GW[78] GW[79] GW[80]
+ GW[81] GW[82] GW[83] GW[84] GW[85] GW[86] GW[87] GW[88] GW[89] GW[90] GW[91]
+ GW[92] GW[93] GW[94] GW[95] GW[96] GW[97] GW[98] GW[99] GW[100] GW[101]
+ GW[102] GW[103] GW[104] GW[105] GW[106] GW[107] GW[108] GW[109] GW[110]
+ GW[111] GW[112] GW[113] GW[114] GW[115] GW[116] GW[117] GW[118] GW[119]
+ GW[120] GW[121] GW[122] GW[123] GW[124] GW[125] GW[126] GW[127] GWB[69]
+ GWB[70] GWB[71] GWB[72] GWB[73] GWB[74] GWB[75] GWB[76] GWB[77] GWB[78]
+ GWB[79] GWB[80] GWB[81] GWB[82] GWB[83] GWB[84] GWB[85] GWB[86] GWB[87]
+ GWB[88] GWB[89] GWB[90] GWB[91] GWB[92] GWB[93] GWB[94] GWB[95] GWB[96]
+ GWB[97] GWB[98] GWB[99] GWB[100] GWB[101] GWB[102] GWB[103] GWB[104] GWB[105]
+ GWB[106] GWB[107] GWB[108] GWB[109] GWB[110] GWB[111] GWB[112] GWB[113]
+ GWB[114] GWB[115] GWB[116] GWB[117] GWB[118] GWB[119] GWB[120] GWB[121]
+ GWB[122] GWB[123] GWB[124] GWB[125] GWB[126] GWB[127] PHASESEL_R QA[69] QA[70]
+ QA[71] QA[72] QA[73] QA[74] QA[75] QA[76] QA[77] QA[78] QA[79] QA[80] QA[81]
+ QA[82] QA[83] QA[84] QA[85] QA[86] QA[87] QA[88] QA[89] QA[90] QA[91] QA[92]
+ QA[93] QA[94] QA[95] QA[96] QA[97] QA[98] QA[99] QA[100] QA[101] QA[102]
+ QA[103] QA[104] QA[105] QA[106] QA[107] QA[108] QA[109] QA[110] QA[111]
+ QA[112] QA[113] QA[114] QA[115] QA[116] QA[117] QA[118] QA[119] QA[120]
+ QA[121] QA[122] QA[123] QA[124] QA[125] QA[126] QA[127] QB[69] QB[70] QB[71]
+ QB[72] QB[73] QB[74] QB[75] QB[76] QB[77] QB[78] QB[79] QB[80] QB[81] QB[82]
+ QB[83] QB[84] QB[85] QB[86] QB[87] QB[88] QB[89] QB[90] QB[91] QB[92] QB[93]
+ QB[94] QB[95] QB[96] QB[97] QB[98] QB[99] QB[100] QB[101] QB[102] QB[103]
+ QB[104] QB[105] QB[106] QB[107] QB[108] QB[109] QB[110] QB[111] QB[112]
+ QB[113] QB[114] QB[115] QB[116] QB[117] QB[118] QB[119] QB[120] QB[121]
+ QB[122] QB[123] QB[124] QB[125] QB[126] QB[127] QLATCH_AB_R QLATCH_BB_R
+ RSC_TRK_W VDD VSS VLO WLP_SAEB SDBM200W80_MIO_R
XCNT_CORE_IO_M4 VLO AWT2 BLTRKWLDRV CEBA CEBB CKD CLK DCLKA DCLK_L DCLK_R
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X3[0] DEC_X3[1] DEC_X3[2]
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2]
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PHASESEL_L PHASESEL_R PTSEL[0]
+ PTSEL[1] QLATCH_AB_L QLATCH_AB_R QLATCH_BB_L QLATCH_BB_R RSC_TRK_W RTSEL[0]
+ RTSEL[1] VLO VLO TRKBL VDD VHI VLO VSS WEBA WEBB WLP_SAE WLP_SAEB WLP_SAE_TK
+ WTSEL[0] WTSEL[1] AA[2] AA[3] AA[4] AA[5] AA[6] AA[7] VLO AA[8] VLO VLO AB[2]
+ AB[3] AB[4] AB[5] AB[6] AB[7] VLO AB[8] VLO VLO AA[0] AA[1] AB[0] AB[1] VLO
+ VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO
+ DA[59] DA[60] DA[61] DA[62] DA[63] DA[64] DA[65] DA[66] DA[67] DA[68] DB[59]
+ DB[60] DB[61] DB[62] DB[63] DB[64] DB[65] DB[66] DB[67] DB[68] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBL[64] GBL[65] GBL[66] GBL[67] GBL[68] GBLB[59]
+ GBLB[60] GBLB[61] GBLB[62] GBLB[63] GBLB[64] GBLB[65] GBLB[66] GBLB[67]
+ GBLB[68] GW[59] GW[60] GW[61] GW[62] GW[63] GW[64] GW[65] GW[66] GW[67] GW[68]
+ GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] GWB[64] GWB[65] GWB[66] GWB[67]
+ GWB[68] QA[59] QA[60] QA[61] QA[62] QA[63] QA[64] QA[65] QA[66] QA[67] QA[68]
+ QB[59] QB[60] QB[61] QB[62] QB[63] QB[64] QB[65] QB[66] QB[67] QB[68]
+ SDBM200W80_CNT_CORE_IO
XTOPEDGE VDD VSS WLP_SAE WLP_SAE_TK SDBM200W80_TOP_EDGE
XD_WEBA WEBA VSS SDBM200W80_DIO
XD_WEBB WEBB VSS SDBM200W80_DIO
XD_CEBA CEBA VSS SDBM200W80_DIO
XD_CEBB CEBB VSS SDBM200W80_DIO
XD_WTESL_1 WTSEL[1] VSS SDBM200W80_DIO
XD_WTESL_0 WTSEL[0] VSS SDBM200W80_DIO
XD_RTESL_1 RTSEL[1] VSS SDBM200W80_DIO
XD_RTESL_0 RTSEL[0] VSS SDBM200W80_DIO
XD_PTESL_1 PTSEL[1] VSS SDBM200W80_DIO
XD_PTESL_0 PTSEL[0] VSS SDBM200W80_DIO
XD_CLK CLK VSS SDBM200W80_DIO
XD_AA0 AA[0] VSS SDBM200W80_DIO
XD_AA1 AA[1] VSS SDBM200W80_DIO
XD_AA2 AA[2] VSS SDBM200W80_DIO
XD_AA3 AA[3] VSS SDBM200W80_DIO
XD_AA4 AA[4] VSS SDBM200W80_DIO
XD_AA5 AA[5] VSS SDBM200W80_DIO
XD_AA6 AA[6] VSS SDBM200W80_DIO
XD_AA7 AA[7] VSS SDBM200W80_DIO
XD_AA8 AA[8] VSS SDBM200W80_DIO
XD_AB0 AB[0] VSS SDBM200W80_DIO
XD_AB1 AB[1] VSS SDBM200W80_DIO
XD_AB2 AB[2] VSS SDBM200W80_DIO
XD_AB3 AB[3] VSS SDBM200W80_DIO
XD_AB4 AB[4] VSS SDBM200W80_DIO
XD_AB5 AB[5] VSS SDBM200W80_DIO
XD_AB6 AB[6] VSS SDBM200W80_DIO
XD_AB7 AB[7] VSS SDBM200W80_DIO
XD_AB8 AB[8] VSS SDBM200W80_DIO
XD_DA0 DA[0] VSS SDBM200W80_DIO
XD_DA1 DA[1] VSS SDBM200W80_DIO
XD_DA2 DA[2] VSS SDBM200W80_DIO
XD_DA3 DA[3] VSS SDBM200W80_DIO
XD_DA4 DA[4] VSS SDBM200W80_DIO
XD_DA5 DA[5] VSS SDBM200W80_DIO
XD_DA6 DA[6] VSS SDBM200W80_DIO
XD_DA7 DA[7] VSS SDBM200W80_DIO
XD_DA8 DA[8] VSS SDBM200W80_DIO
XD_DA9 DA[9] VSS SDBM200W80_DIO
XD_DA10 DA[10] VSS SDBM200W80_DIO
XD_DA11 DA[11] VSS SDBM200W80_DIO
XD_DA12 DA[12] VSS SDBM200W80_DIO
XD_DA13 DA[13] VSS SDBM200W80_DIO
XD_DA14 DA[14] VSS SDBM200W80_DIO
XD_DA15 DA[15] VSS SDBM200W80_DIO
XD_DA16 DA[16] VSS SDBM200W80_DIO
XD_DA17 DA[17] VSS SDBM200W80_DIO
XD_DA18 DA[18] VSS SDBM200W80_DIO
XD_DA19 DA[19] VSS SDBM200W80_DIO
XD_DA20 DA[20] VSS SDBM200W80_DIO
XD_DA21 DA[21] VSS SDBM200W80_DIO
XD_DA22 DA[22] VSS SDBM200W80_DIO
XD_DA23 DA[23] VSS SDBM200W80_DIO
XD_DA24 DA[24] VSS SDBM200W80_DIO
XD_DA25 DA[25] VSS SDBM200W80_DIO
XD_DA26 DA[26] VSS SDBM200W80_DIO
XD_DA27 DA[27] VSS SDBM200W80_DIO
XD_DA28 DA[28] VSS SDBM200W80_DIO
XD_DA29 DA[29] VSS SDBM200W80_DIO
XD_DA30 DA[30] VSS SDBM200W80_DIO
XD_DA31 DA[31] VSS SDBM200W80_DIO
XD_DA32 DA[32] VSS SDBM200W80_DIO
XD_DA33 DA[33] VSS SDBM200W80_DIO
XD_DA34 DA[34] VSS SDBM200W80_DIO
XD_DA35 DA[35] VSS SDBM200W80_DIO
XD_DA36 DA[36] VSS SDBM200W80_DIO
XD_DA37 DA[37] VSS SDBM200W80_DIO
XD_DA38 DA[38] VSS SDBM200W80_DIO
XD_DA39 DA[39] VSS SDBM200W80_DIO
XD_DA40 DA[40] VSS SDBM200W80_DIO
XD_DA41 DA[41] VSS SDBM200W80_DIO
XD_DA42 DA[42] VSS SDBM200W80_DIO
XD_DA43 DA[43] VSS SDBM200W80_DIO
XD_DA44 DA[44] VSS SDBM200W80_DIO
XD_DA45 DA[45] VSS SDBM200W80_DIO
XD_DA46 DA[46] VSS SDBM200W80_DIO
XD_DA47 DA[47] VSS SDBM200W80_DIO
XD_DA48 DA[48] VSS SDBM200W80_DIO
XD_DA49 DA[49] VSS SDBM200W80_DIO
XD_DA50 DA[50] VSS SDBM200W80_DIO
XD_DA51 DA[51] VSS SDBM200W80_DIO
XD_DA52 DA[52] VSS SDBM200W80_DIO
XD_DA53 DA[53] VSS SDBM200W80_DIO
XD_DA54 DA[54] VSS SDBM200W80_DIO
XD_DA55 DA[55] VSS SDBM200W80_DIO
XD_DA56 DA[56] VSS SDBM200W80_DIO
XD_DA57 DA[57] VSS SDBM200W80_DIO
XD_DA58 DA[58] VSS SDBM200W80_DIO
XD_DA59 DA[59] VSS SDBM200W80_DIO
XD_DA60 DA[60] VSS SDBM200W80_DIO
XD_DA61 DA[61] VSS SDBM200W80_DIO
XD_DA62 DA[62] VSS SDBM200W80_DIO
XD_DA63 DA[63] VSS SDBM200W80_DIO
XD_DA64 DA[64] VSS SDBM200W80_DIO
XD_DA65 DA[65] VSS SDBM200W80_DIO
XD_DA66 DA[66] VSS SDBM200W80_DIO
XD_DA67 DA[67] VSS SDBM200W80_DIO
XD_DA68 DA[68] VSS SDBM200W80_DIO
XD_DA69 DA[69] VSS SDBM200W80_DIO
XD_DA70 DA[70] VSS SDBM200W80_DIO
XD_DA71 DA[71] VSS SDBM200W80_DIO
XD_DA72 DA[72] VSS SDBM200W80_DIO
XD_DA73 DA[73] VSS SDBM200W80_DIO
XD_DA74 DA[74] VSS SDBM200W80_DIO
XD_DA75 DA[75] VSS SDBM200W80_DIO
XD_DA76 DA[76] VSS SDBM200W80_DIO
XD_DA77 DA[77] VSS SDBM200W80_DIO
XD_DA78 DA[78] VSS SDBM200W80_DIO
XD_DA79 DA[79] VSS SDBM200W80_DIO
XD_DA80 DA[80] VSS SDBM200W80_DIO
XD_DA81 DA[81] VSS SDBM200W80_DIO
XD_DA82 DA[82] VSS SDBM200W80_DIO
XD_DA83 DA[83] VSS SDBM200W80_DIO
XD_DA84 DA[84] VSS SDBM200W80_DIO
XD_DA85 DA[85] VSS SDBM200W80_DIO
XD_DA86 DA[86] VSS SDBM200W80_DIO
XD_DA87 DA[87] VSS SDBM200W80_DIO
XD_DA88 DA[88] VSS SDBM200W80_DIO
XD_DA89 DA[89] VSS SDBM200W80_DIO
XD_DA90 DA[90] VSS SDBM200W80_DIO
XD_DA91 DA[91] VSS SDBM200W80_DIO
XD_DA92 DA[92] VSS SDBM200W80_DIO
XD_DA93 DA[93] VSS SDBM200W80_DIO
XD_DA94 DA[94] VSS SDBM200W80_DIO
XD_DA95 DA[95] VSS SDBM200W80_DIO
XD_DA96 DA[96] VSS SDBM200W80_DIO
XD_DA97 DA[97] VSS SDBM200W80_DIO
XD_DA98 DA[98] VSS SDBM200W80_DIO
XD_DA99 DA[99] VSS SDBM200W80_DIO
XD_DA100 DA[100] VSS SDBM200W80_DIO
XD_DA101 DA[101] VSS SDBM200W80_DIO
XD_DA102 DA[102] VSS SDBM200W80_DIO
XD_DA103 DA[103] VSS SDBM200W80_DIO
XD_DA104 DA[104] VSS SDBM200W80_DIO
XD_DA105 DA[105] VSS SDBM200W80_DIO
XD_DA106 DA[106] VSS SDBM200W80_DIO
XD_DA107 DA[107] VSS SDBM200W80_DIO
XD_DA108 DA[108] VSS SDBM200W80_DIO
XD_DA109 DA[109] VSS SDBM200W80_DIO
XD_DA110 DA[110] VSS SDBM200W80_DIO
XD_DA111 DA[111] VSS SDBM200W80_DIO
XD_DA112 DA[112] VSS SDBM200W80_DIO
XD_DA113 DA[113] VSS SDBM200W80_DIO
XD_DA114 DA[114] VSS SDBM200W80_DIO
XD_DA115 DA[115] VSS SDBM200W80_DIO
XD_DA116 DA[116] VSS SDBM200W80_DIO
XD_DA117 DA[117] VSS SDBM200W80_DIO
XD_DA118 DA[118] VSS SDBM200W80_DIO
XD_DA119 DA[119] VSS SDBM200W80_DIO
XD_DA120 DA[120] VSS SDBM200W80_DIO
XD_DA121 DA[121] VSS SDBM200W80_DIO
XD_DA122 DA[122] VSS SDBM200W80_DIO
XD_DA123 DA[123] VSS SDBM200W80_DIO
XD_DA124 DA[124] VSS SDBM200W80_DIO
XD_DA125 DA[125] VSS SDBM200W80_DIO
XD_DA126 DA[126] VSS SDBM200W80_DIO
XD_DA127 DA[127] VSS SDBM200W80_DIO
XD_DB0 DB[0] VSS SDBM200W80_DIO
XD_DB1 DB[1] VSS SDBM200W80_DIO
XD_DB2 DB[2] VSS SDBM200W80_DIO
XD_DB3 DB[3] VSS SDBM200W80_DIO
XD_DB4 DB[4] VSS SDBM200W80_DIO
XD_DB5 DB[5] VSS SDBM200W80_DIO
XD_DB6 DB[6] VSS SDBM200W80_DIO
XD_DB7 DB[7] VSS SDBM200W80_DIO
XD_DB8 DB[8] VSS SDBM200W80_DIO
XD_DB9 DB[9] VSS SDBM200W80_DIO
XD_DB10 DB[10] VSS SDBM200W80_DIO
XD_DB11 DB[11] VSS SDBM200W80_DIO
XD_DB12 DB[12] VSS SDBM200W80_DIO
XD_DB13 DB[13] VSS SDBM200W80_DIO
XD_DB14 DB[14] VSS SDBM200W80_DIO
XD_DB15 DB[15] VSS SDBM200W80_DIO
XD_DB16 DB[16] VSS SDBM200W80_DIO
XD_DB17 DB[17] VSS SDBM200W80_DIO
XD_DB18 DB[18] VSS SDBM200W80_DIO
XD_DB19 DB[19] VSS SDBM200W80_DIO
XD_DB20 DB[20] VSS SDBM200W80_DIO
XD_DB21 DB[21] VSS SDBM200W80_DIO
XD_DB22 DB[22] VSS SDBM200W80_DIO
XD_DB23 DB[23] VSS SDBM200W80_DIO
XD_DB24 DB[24] VSS SDBM200W80_DIO
XD_DB25 DB[25] VSS SDBM200W80_DIO
XD_DB26 DB[26] VSS SDBM200W80_DIO
XD_DB27 DB[27] VSS SDBM200W80_DIO
XD_DB28 DB[28] VSS SDBM200W80_DIO
XD_DB29 DB[29] VSS SDBM200W80_DIO
XD_DB30 DB[30] VSS SDBM200W80_DIO
XD_DB31 DB[31] VSS SDBM200W80_DIO
XD_DB32 DB[32] VSS SDBM200W80_DIO
XD_DB33 DB[33] VSS SDBM200W80_DIO
XD_DB34 DB[34] VSS SDBM200W80_DIO
XD_DB35 DB[35] VSS SDBM200W80_DIO
XD_DB36 DB[36] VSS SDBM200W80_DIO
XD_DB37 DB[37] VSS SDBM200W80_DIO
XD_DB38 DB[38] VSS SDBM200W80_DIO
XD_DB39 DB[39] VSS SDBM200W80_DIO
XD_DB40 DB[40] VSS SDBM200W80_DIO
XD_DB41 DB[41] VSS SDBM200W80_DIO
XD_DB42 DB[42] VSS SDBM200W80_DIO
XD_DB43 DB[43] VSS SDBM200W80_DIO
XD_DB44 DB[44] VSS SDBM200W80_DIO
XD_DB45 DB[45] VSS SDBM200W80_DIO
XD_DB46 DB[46] VSS SDBM200W80_DIO
XD_DB47 DB[47] VSS SDBM200W80_DIO
XD_DB48 DB[48] VSS SDBM200W80_DIO
XD_DB49 DB[49] VSS SDBM200W80_DIO
XD_DB50 DB[50] VSS SDBM200W80_DIO
XD_DB51 DB[51] VSS SDBM200W80_DIO
XD_DB52 DB[52] VSS SDBM200W80_DIO
XD_DB53 DB[53] VSS SDBM200W80_DIO
XD_DB54 DB[54] VSS SDBM200W80_DIO
XD_DB55 DB[55] VSS SDBM200W80_DIO
XD_DB56 DB[56] VSS SDBM200W80_DIO
XD_DB57 DB[57] VSS SDBM200W80_DIO
XD_DB58 DB[58] VSS SDBM200W80_DIO
XD_DB59 DB[59] VSS SDBM200W80_DIO
XD_DB60 DB[60] VSS SDBM200W80_DIO
XD_DB61 DB[61] VSS SDBM200W80_DIO
XD_DB62 DB[62] VSS SDBM200W80_DIO
XD_DB63 DB[63] VSS SDBM200W80_DIO
XD_DB64 DB[64] VSS SDBM200W80_DIO
XD_DB65 DB[65] VSS SDBM200W80_DIO
XD_DB66 DB[66] VSS SDBM200W80_DIO
XD_DB67 DB[67] VSS SDBM200W80_DIO
XD_DB68 DB[68] VSS SDBM200W80_DIO
XD_DB69 DB[69] VSS SDBM200W80_DIO
XD_DB70 DB[70] VSS SDBM200W80_DIO
XD_DB71 DB[71] VSS SDBM200W80_DIO
XD_DB72 DB[72] VSS SDBM200W80_DIO
XD_DB73 DB[73] VSS SDBM200W80_DIO
XD_DB74 DB[74] VSS SDBM200W80_DIO
XD_DB75 DB[75] VSS SDBM200W80_DIO
XD_DB76 DB[76] VSS SDBM200W80_DIO
XD_DB77 DB[77] VSS SDBM200W80_DIO
XD_DB78 DB[78] VSS SDBM200W80_DIO
XD_DB79 DB[79] VSS SDBM200W80_DIO
XD_DB80 DB[80] VSS SDBM200W80_DIO
XD_DB81 DB[81] VSS SDBM200W80_DIO
XD_DB82 DB[82] VSS SDBM200W80_DIO
XD_DB83 DB[83] VSS SDBM200W80_DIO
XD_DB84 DB[84] VSS SDBM200W80_DIO
XD_DB85 DB[85] VSS SDBM200W80_DIO
XD_DB86 DB[86] VSS SDBM200W80_DIO
XD_DB87 DB[87] VSS SDBM200W80_DIO
XD_DB88 DB[88] VSS SDBM200W80_DIO
XD_DB89 DB[89] VSS SDBM200W80_DIO
XD_DB90 DB[90] VSS SDBM200W80_DIO
XD_DB91 DB[91] VSS SDBM200W80_DIO
XD_DB92 DB[92] VSS SDBM200W80_DIO
XD_DB93 DB[93] VSS SDBM200W80_DIO
XD_DB94 DB[94] VSS SDBM200W80_DIO
XD_DB95 DB[95] VSS SDBM200W80_DIO
XD_DB96 DB[96] VSS SDBM200W80_DIO
XD_DB97 DB[97] VSS SDBM200W80_DIO
XD_DB98 DB[98] VSS SDBM200W80_DIO
XD_DB99 DB[99] VSS SDBM200W80_DIO
XD_DB100 DB[100] VSS SDBM200W80_DIO
XD_DB101 DB[101] VSS SDBM200W80_DIO
XD_DB102 DB[102] VSS SDBM200W80_DIO
XD_DB103 DB[103] VSS SDBM200W80_DIO
XD_DB104 DB[104] VSS SDBM200W80_DIO
XD_DB105 DB[105] VSS SDBM200W80_DIO
XD_DB106 DB[106] VSS SDBM200W80_DIO
XD_DB107 DB[107] VSS SDBM200W80_DIO
XD_DB108 DB[108] VSS SDBM200W80_DIO
XD_DB109 DB[109] VSS SDBM200W80_DIO
XD_DB110 DB[110] VSS SDBM200W80_DIO
XD_DB111 DB[111] VSS SDBM200W80_DIO
XD_DB112 DB[112] VSS SDBM200W80_DIO
XD_DB113 DB[113] VSS SDBM200W80_DIO
XD_DB114 DB[114] VSS SDBM200W80_DIO
XD_DB115 DB[115] VSS SDBM200W80_DIO
XD_DB116 DB[116] VSS SDBM200W80_DIO
XD_DB117 DB[117] VSS SDBM200W80_DIO
XD_DB118 DB[118] VSS SDBM200W80_DIO
XD_DB119 DB[119] VSS SDBM200W80_DIO
XD_DB120 DB[120] VSS SDBM200W80_DIO
XD_DB121 DB[121] VSS SDBM200W80_DIO
XD_DB122 DB[122] VSS SDBM200W80_DIO
XD_DB123 DB[123] VSS SDBM200W80_DIO
XD_DB124 DB[124] VSS SDBM200W80_DIO
XD_DB125 DB[125] VSS SDBM200W80_DIO
XD_DB126 DB[126] VSS SDBM200W80_DIO
XD_DB127 DB[127] VSS SDBM200W80_DIO
.ENDS

