# Created by MC2 : Version 2012.02.00.d on 2024/01/10, 17:24:41

#*********************************************************************************************************************/
# Software       : TSMC MEMORY COMPILER tsn28hpcpuhddpsram_2012.02.00.d.170a						*/
# Technology     : TSMC 28nm CMOS LOGIC High Performance Compact Mobile 1P10M HKMG CU_ELK 0.9V				*/
# Memory Type    : TSMC 28nm High Performance Compact Mobile Ultra High Density Dual Port SRAM with d127 bit cell SVT Periphery */
# Library Name   : tsdn28hpcpuhdb512x128m4m (user specify : TSDN28HPCPUHDB512X128M4M)				*/
# Library Version: 170a												*/
# Generated Time : 2024/01/10, 17:23:40										*/
#*********************************************************************************************************************/
#															*/
# STATEMENT OF USE													*/
#															*/
# This information contains confidential and proprietary information of TSMC.					*/
# No part of this information may be reproduced, transmitted, transcribed,						*/
# stored in a retrieval system, or translated into any human or computer						*/
# language, in any form or by any means, electronic, mechanical, magnetic,						*/
# optical, chemical, manual, or otherwise, without the prior written permission					*/
# of TSMC. This information was prepared for informational purpose and is for					*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the					*/
# information at any time and without notice.									*/
#															*/
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TSDN28HPCPUHDB512X128M4M
	CLASS BLOCK ;
	FOREIGN TSDN28HPCPUHDB512X128M4M 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 80.475 BY 317.690 ;
	SYMMETRY X Y ;
	PIN AA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 159.485 80.475 159.635 ;
			LAYER M1 ;
			RECT 80.295 159.485 80.475 159.635 ;
			LAYER M2 ;
			RECT 80.295 159.485 80.475 159.635 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[0]

	PIN AA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 162.035 80.475 162.185 ;
			LAYER M3 ;
			RECT 80.295 162.035 80.475 162.185 ;
			LAYER M1 ;
			RECT 80.295 162.035 80.475 162.185 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[1]

	PIN AA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 151.935 80.475 152.085 ;
			LAYER M2 ;
			RECT 80.295 151.935 80.475 152.085 ;
			LAYER M3 ;
			RECT 80.295 151.935 80.475 152.085 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[2]

	PIN AA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 153.385 80.475 153.535 ;
			LAYER M1 ;
			RECT 80.295 153.385 80.475 153.535 ;
			LAYER M3 ;
			RECT 80.295 153.385 80.475 153.535 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[3]

	PIN AA[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 153.745 80.475 153.895 ;
			LAYER M1 ;
			RECT 80.295 153.745 80.475 153.895 ;
			LAYER M2 ;
			RECT 80.295 153.745 80.475 153.895 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[4]

	PIN AA[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 154.785 80.475 154.935 ;
			LAYER M1 ;
			RECT 80.295 154.785 80.475 154.935 ;
			LAYER M2 ;
			RECT 80.295 154.785 80.475 154.935 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[5]

	PIN AA[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 156.700 80.475 156.850 ;
			LAYER M2 ;
			RECT 80.295 156.700 80.475 156.850 ;
			LAYER M1 ;
			RECT 80.295 156.700 80.475 156.850 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[6]

	PIN AA[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 157.255 80.475 157.405 ;
			LAYER M3 ;
			RECT 80.295 157.255 80.475 157.405 ;
			LAYER M1 ;
			RECT 80.295 157.255 80.475 157.405 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[7]

	PIN AA[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 163.025 80.475 163.175 ;
			LAYER M3 ;
			RECT 80.295 163.025 80.475 163.175 ;
			LAYER M1 ;
			RECT 80.295 163.025 80.475 163.175 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[8]

	PIN AB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 159.815 80.475 159.965 ;
			LAYER M3 ;
			RECT 80.295 159.815 80.475 159.965 ;
			LAYER M1 ;
			RECT 80.295 159.815 80.475 159.965 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[0]

	PIN AB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 161.705 80.475 161.855 ;
			LAYER M2 ;
			RECT 80.295 161.705 80.475 161.855 ;
			LAYER M3 ;
			RECT 80.295 161.705 80.475 161.855 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[1]

	PIN AB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 152.265 80.475 152.415 ;
			LAYER M2 ;
			RECT 80.295 152.265 80.475 152.415 ;
			LAYER M1 ;
			RECT 80.295 152.265 80.475 152.415 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[2]

	PIN AB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 153.055 80.475 153.205 ;
			LAYER M3 ;
			RECT 80.295 153.055 80.475 153.205 ;
			LAYER M1 ;
			RECT 80.295 153.055 80.475 153.205 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[3]

	PIN AB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 154.075 80.475 154.225 ;
			LAYER M1 ;
			RECT 80.295 154.075 80.475 154.225 ;
			LAYER M3 ;
			RECT 80.295 154.075 80.475 154.225 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[4]

	PIN AB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 155.945 80.475 156.095 ;
			LAYER M1 ;
			RECT 80.295 155.945 80.475 156.095 ;
			LAYER M3 ;
			RECT 80.295 155.945 80.475 156.095 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[5]

	PIN AB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 156.370 80.475 156.520 ;
			LAYER M1 ;
			RECT 80.295 156.370 80.475 156.520 ;
			LAYER M2 ;
			RECT 80.295 156.370 80.475 156.520 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[6]

	PIN AB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 157.585 80.475 157.735 ;
			LAYER M2 ;
			RECT 80.295 157.585 80.475 157.735 ;
			LAYER M3 ;
			RECT 80.295 157.585 80.475 157.735 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[7]

	PIN AB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 163.355 80.475 163.505 ;
			LAYER M3 ;
			RECT 80.295 163.355 80.475 163.505 ;
			LAYER M2 ;
			RECT 80.295 163.355 80.475 163.505 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[8]

	PIN CEBA
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 166.620 80.475 166.770 ;
			LAYER M2 ;
			RECT 80.295 166.620 80.475 166.770 ;
			LAYER M1 ;
			RECT 80.295 166.620 80.475 166.770 ;
		END
		ANTENNAGATEAREA 0.068100 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.266600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.847400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.223400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.068100 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.577800 LAYER M2 ;
		ANTENNAMAXAREACAR 10.714500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.318800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.068100 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.261500 LAYER M3 ;
		ANTENNAMAXAREACAR 12.155100 LAYER M3 ;
	END CEBA

	PIN CEBB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 166.950 80.475 167.100 ;
			LAYER M2 ;
			RECT 80.295 166.950 80.475 167.100 ;
			LAYER M3 ;
			RECT 80.295 166.950 80.475 167.100 ;
		END
		ANTENNAGATEAREA 0.029100 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.342200 LAYER M1 ;
		ANTENNAMAXAREACAR 10.096200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.223400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.029100 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.644400 LAYER M2 ;
		ANTENNAMAXAREACAR 32.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.446700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.029100 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 33.167500 LAYER M3 ;
	END CEBB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 164.640 80.475 164.790 ;
			LAYER M1 ;
			RECT 80.295 164.640 80.475 164.790 ;
			LAYER M2 ;
			RECT 80.295 164.640 80.475 164.790 ;
		END
		ANTENNAGATEAREA 0.394500 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.757100 LAYER M1 ;
		ANTENNAMAXAREACAR 3.389600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.656600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.394500 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.828600 LAYER M2 ;
		ANTENNAMAXAREACAR 8.667400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.313100 LAYER VIA2 ;
		ANTENNAGATEAREA 0.394500 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.952600 LAYER M3 ;
		ANTENNAMAXAREACAR 11.082000 LAYER M3 ;
	END CLK

	PIN DA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 2.855 80.475 3.005 ;
			LAYER M2 ;
			RECT 80.295 2.855 80.475 3.005 ;
			LAYER M1 ;
			RECT 80.295 2.855 80.475 3.005 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[0]

	PIN DA[100]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 253.375 80.475 253.525 ;
			LAYER M3 ;
			RECT 80.295 253.375 80.475 253.525 ;
			LAYER M1 ;
			RECT 80.295 253.375 80.475 253.525 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[100]

	PIN DA[101]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 255.695 80.475 255.845 ;
			LAYER M1 ;
			RECT 80.295 255.695 80.475 255.845 ;
			LAYER M3 ;
			RECT 80.295 255.695 80.475 255.845 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[101]

	PIN DA[102]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 258.015 80.475 258.165 ;
			LAYER M3 ;
			RECT 80.295 258.015 80.475 258.165 ;
			LAYER M2 ;
			RECT 80.295 258.015 80.475 258.165 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[102]

	PIN DA[103]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 260.335 80.475 260.485 ;
			LAYER M1 ;
			RECT 80.295 260.335 80.475 260.485 ;
			LAYER M2 ;
			RECT 80.295 260.335 80.475 260.485 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[103]

	PIN DA[104]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 262.655 80.475 262.805 ;
			LAYER M1 ;
			RECT 80.295 262.655 80.475 262.805 ;
			LAYER M3 ;
			RECT 80.295 262.655 80.475 262.805 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[104]

	PIN DA[105]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 264.975 80.475 265.125 ;
			LAYER M3 ;
			RECT 80.295 264.975 80.475 265.125 ;
			LAYER M2 ;
			RECT 80.295 264.975 80.475 265.125 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[105]

	PIN DA[106]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 267.295 80.475 267.445 ;
			LAYER M3 ;
			RECT 80.295 267.295 80.475 267.445 ;
			LAYER M2 ;
			RECT 80.295 267.295 80.475 267.445 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[106]

	PIN DA[107]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 269.615 80.475 269.765 ;
			LAYER M3 ;
			RECT 80.295 269.615 80.475 269.765 ;
			LAYER M1 ;
			RECT 80.295 269.615 80.475 269.765 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[107]

	PIN DA[108]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 271.935 80.475 272.085 ;
			LAYER M1 ;
			RECT 80.295 271.935 80.475 272.085 ;
			LAYER M3 ;
			RECT 80.295 271.935 80.475 272.085 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[108]

	PIN DA[109]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 274.255 80.475 274.405 ;
			LAYER M2 ;
			RECT 80.295 274.255 80.475 274.405 ;
			LAYER M3 ;
			RECT 80.295 274.255 80.475 274.405 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[109]

	PIN DA[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 26.055 80.475 26.205 ;
			LAYER M3 ;
			RECT 80.295 26.055 80.475 26.205 ;
			LAYER M2 ;
			RECT 80.295 26.055 80.475 26.205 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[10]

	PIN DA[110]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 276.575 80.475 276.725 ;
			LAYER M3 ;
			RECT 80.295 276.575 80.475 276.725 ;
			LAYER M2 ;
			RECT 80.295 276.575 80.475 276.725 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[110]

	PIN DA[111]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 278.895 80.475 279.045 ;
			LAYER M2 ;
			RECT 80.295 278.895 80.475 279.045 ;
			LAYER M3 ;
			RECT 80.295 278.895 80.475 279.045 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[111]

	PIN DA[112]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 281.215 80.475 281.365 ;
			LAYER M1 ;
			RECT 80.295 281.215 80.475 281.365 ;
			LAYER M2 ;
			RECT 80.295 281.215 80.475 281.365 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[112]

	PIN DA[113]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 283.535 80.475 283.685 ;
			LAYER M2 ;
			RECT 80.295 283.535 80.475 283.685 ;
			LAYER M3 ;
			RECT 80.295 283.535 80.475 283.685 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[113]

	PIN DA[114]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 285.855 80.475 286.005 ;
			LAYER M2 ;
			RECT 80.295 285.855 80.475 286.005 ;
			LAYER M1 ;
			RECT 80.295 285.855 80.475 286.005 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[114]

	PIN DA[115]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 288.175 80.475 288.325 ;
			LAYER M2 ;
			RECT 80.295 288.175 80.475 288.325 ;
			LAYER M1 ;
			RECT 80.295 288.175 80.475 288.325 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[115]

	PIN DA[116]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 290.495 80.475 290.645 ;
			LAYER M3 ;
			RECT 80.295 290.495 80.475 290.645 ;
			LAYER M1 ;
			RECT 80.295 290.495 80.475 290.645 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[116]

	PIN DA[117]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 292.815 80.475 292.965 ;
			LAYER M3 ;
			RECT 80.295 292.815 80.475 292.965 ;
			LAYER M1 ;
			RECT 80.295 292.815 80.475 292.965 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[117]

	PIN DA[118]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 295.135 80.475 295.285 ;
			LAYER M2 ;
			RECT 80.295 295.135 80.475 295.285 ;
			LAYER M3 ;
			RECT 80.295 295.135 80.475 295.285 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[118]

	PIN DA[119]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 297.455 80.475 297.605 ;
			LAYER M2 ;
			RECT 80.295 297.455 80.475 297.605 ;
			LAYER M1 ;
			RECT 80.295 297.455 80.475 297.605 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[119]

	PIN DA[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 28.375 80.475 28.525 ;
			LAYER M2 ;
			RECT 80.295 28.375 80.475 28.525 ;
			LAYER M1 ;
			RECT 80.295 28.375 80.475 28.525 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[11]

	PIN DA[120]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 299.775 80.475 299.925 ;
			LAYER M3 ;
			RECT 80.295 299.775 80.475 299.925 ;
			LAYER M1 ;
			RECT 80.295 299.775 80.475 299.925 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[120]

	PIN DA[121]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 302.095 80.475 302.245 ;
			LAYER M3 ;
			RECT 80.295 302.095 80.475 302.245 ;
			LAYER M1 ;
			RECT 80.295 302.095 80.475 302.245 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[121]

	PIN DA[122]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 304.415 80.475 304.565 ;
			LAYER M2 ;
			RECT 80.295 304.415 80.475 304.565 ;
			LAYER M1 ;
			RECT 80.295 304.415 80.475 304.565 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[122]

	PIN DA[123]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 306.735 80.475 306.885 ;
			LAYER M3 ;
			RECT 80.295 306.735 80.475 306.885 ;
			LAYER M2 ;
			RECT 80.295 306.735 80.475 306.885 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[123]

	PIN DA[124]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 309.055 80.475 309.205 ;
			LAYER M2 ;
			RECT 80.295 309.055 80.475 309.205 ;
			LAYER M3 ;
			RECT 80.295 309.055 80.475 309.205 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[124]

	PIN DA[125]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 311.375 80.475 311.525 ;
			LAYER M1 ;
			RECT 80.295 311.375 80.475 311.525 ;
			LAYER M2 ;
			RECT 80.295 311.375 80.475 311.525 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[125]

	PIN DA[126]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 313.695 80.475 313.845 ;
			LAYER M1 ;
			RECT 80.295 313.695 80.475 313.845 ;
			LAYER M3 ;
			RECT 80.295 313.695 80.475 313.845 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[126]

	PIN DA[127]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 316.015 80.475 316.165 ;
			LAYER M1 ;
			RECT 80.295 316.015 80.475 316.165 ;
			LAYER M3 ;
			RECT 80.295 316.015 80.475 316.165 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[127]

	PIN DA[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 30.695 80.475 30.845 ;
			LAYER M1 ;
			RECT 80.295 30.695 80.475 30.845 ;
			LAYER M2 ;
			RECT 80.295 30.695 80.475 30.845 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[12]

	PIN DA[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 33.015 80.475 33.165 ;
			LAYER M1 ;
			RECT 80.295 33.015 80.475 33.165 ;
			LAYER M2 ;
			RECT 80.295 33.015 80.475 33.165 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[13]

	PIN DA[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 35.335 80.475 35.485 ;
			LAYER M1 ;
			RECT 80.295 35.335 80.475 35.485 ;
			LAYER M2 ;
			RECT 80.295 35.335 80.475 35.485 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[14]

	PIN DA[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 37.655 80.475 37.805 ;
			LAYER M1 ;
			RECT 80.295 37.655 80.475 37.805 ;
			LAYER M2 ;
			RECT 80.295 37.655 80.475 37.805 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[15]

	PIN DA[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 39.975 80.475 40.125 ;
			LAYER M3 ;
			RECT 80.295 39.975 80.475 40.125 ;
			LAYER M2 ;
			RECT 80.295 39.975 80.475 40.125 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[16]

	PIN DA[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 42.295 80.475 42.445 ;
			LAYER M1 ;
			RECT 80.295 42.295 80.475 42.445 ;
			LAYER M3 ;
			RECT 80.295 42.295 80.475 42.445 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[17]

	PIN DA[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 44.615 80.475 44.765 ;
			LAYER M3 ;
			RECT 80.295 44.615 80.475 44.765 ;
			LAYER M2 ;
			RECT 80.295 44.615 80.475 44.765 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[18]

	PIN DA[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 46.935 80.475 47.085 ;
			LAYER M2 ;
			RECT 80.295 46.935 80.475 47.085 ;
			LAYER M3 ;
			RECT 80.295 46.935 80.475 47.085 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[19]

	PIN DA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 5.175 80.475 5.325 ;
			LAYER M1 ;
			RECT 80.295 5.175 80.475 5.325 ;
			LAYER M2 ;
			RECT 80.295 5.175 80.475 5.325 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[1]

	PIN DA[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 49.255 80.475 49.405 ;
			LAYER M3 ;
			RECT 80.295 49.255 80.475 49.405 ;
			LAYER M1 ;
			RECT 80.295 49.255 80.475 49.405 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[20]

	PIN DA[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 51.575 80.475 51.725 ;
			LAYER M1 ;
			RECT 80.295 51.575 80.475 51.725 ;
			LAYER M3 ;
			RECT 80.295 51.575 80.475 51.725 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[21]

	PIN DA[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 53.895 80.475 54.045 ;
			LAYER M3 ;
			RECT 80.295 53.895 80.475 54.045 ;
			LAYER M1 ;
			RECT 80.295 53.895 80.475 54.045 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[22]

	PIN DA[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 56.215 80.475 56.365 ;
			LAYER M3 ;
			RECT 80.295 56.215 80.475 56.365 ;
			LAYER M2 ;
			RECT 80.295 56.215 80.475 56.365 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[23]

	PIN DA[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 58.535 80.475 58.685 ;
			LAYER M1 ;
			RECT 80.295 58.535 80.475 58.685 ;
			LAYER M3 ;
			RECT 80.295 58.535 80.475 58.685 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[24]

	PIN DA[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 60.855 80.475 61.005 ;
			LAYER M1 ;
			RECT 80.295 60.855 80.475 61.005 ;
			LAYER M3 ;
			RECT 80.295 60.855 80.475 61.005 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[25]

	PIN DA[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 63.175 80.475 63.325 ;
			LAYER M1 ;
			RECT 80.295 63.175 80.475 63.325 ;
			LAYER M3 ;
			RECT 80.295 63.175 80.475 63.325 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[26]

	PIN DA[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 65.495 80.475 65.645 ;
			LAYER M2 ;
			RECT 80.295 65.495 80.475 65.645 ;
			LAYER M1 ;
			RECT 80.295 65.495 80.475 65.645 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[27]

	PIN DA[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 67.815 80.475 67.965 ;
			LAYER M1 ;
			RECT 80.295 67.815 80.475 67.965 ;
			LAYER M2 ;
			RECT 80.295 67.815 80.475 67.965 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[28]

	PIN DA[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 70.135 80.475 70.285 ;
			LAYER M3 ;
			RECT 80.295 70.135 80.475 70.285 ;
			LAYER M1 ;
			RECT 80.295 70.135 80.475 70.285 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[29]

	PIN DA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 7.495 80.475 7.645 ;
			LAYER M1 ;
			RECT 80.295 7.495 80.475 7.645 ;
			LAYER M2 ;
			RECT 80.295 7.495 80.475 7.645 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[2]

	PIN DA[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 72.455 80.475 72.605 ;
			LAYER M1 ;
			RECT 80.295 72.455 80.475 72.605 ;
			LAYER M3 ;
			RECT 80.295 72.455 80.475 72.605 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[30]

	PIN DA[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 74.775 80.475 74.925 ;
			LAYER M2 ;
			RECT 80.295 74.775 80.475 74.925 ;
			LAYER M3 ;
			RECT 80.295 74.775 80.475 74.925 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[31]

	PIN DA[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 77.095 80.475 77.245 ;
			LAYER M2 ;
			RECT 80.295 77.095 80.475 77.245 ;
			LAYER M3 ;
			RECT 80.295 77.095 80.475 77.245 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[32]

	PIN DA[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 79.415 80.475 79.565 ;
			LAYER M3 ;
			RECT 80.295 79.415 80.475 79.565 ;
			LAYER M1 ;
			RECT 80.295 79.415 80.475 79.565 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[33]

	PIN DA[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 81.735 80.475 81.885 ;
			LAYER M2 ;
			RECT 80.295 81.735 80.475 81.885 ;
			LAYER M3 ;
			RECT 80.295 81.735 80.475 81.885 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[34]

	PIN DA[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 84.055 80.475 84.205 ;
			LAYER M2 ;
			RECT 80.295 84.055 80.475 84.205 ;
			LAYER M3 ;
			RECT 80.295 84.055 80.475 84.205 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[35]

	PIN DA[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 86.375 80.475 86.525 ;
			LAYER M2 ;
			RECT 80.295 86.375 80.475 86.525 ;
			LAYER M1 ;
			RECT 80.295 86.375 80.475 86.525 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[36]

	PIN DA[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 88.695 80.475 88.845 ;
			LAYER M2 ;
			RECT 80.295 88.695 80.475 88.845 ;
			LAYER M3 ;
			RECT 80.295 88.695 80.475 88.845 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[37]

	PIN DA[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 91.015 80.475 91.165 ;
			LAYER M2 ;
			RECT 80.295 91.015 80.475 91.165 ;
			LAYER M3 ;
			RECT 80.295 91.015 80.475 91.165 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[38]

	PIN DA[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 93.335 80.475 93.485 ;
			LAYER M2 ;
			RECT 80.295 93.335 80.475 93.485 ;
			LAYER M3 ;
			RECT 80.295 93.335 80.475 93.485 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[39]

	PIN DA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 9.815 80.475 9.965 ;
			LAYER M2 ;
			RECT 80.295 9.815 80.475 9.965 ;
			LAYER M3 ;
			RECT 80.295 9.815 80.475 9.965 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[3]

	PIN DA[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 95.655 80.475 95.805 ;
			LAYER M2 ;
			RECT 80.295 95.655 80.475 95.805 ;
			LAYER M1 ;
			RECT 80.295 95.655 80.475 95.805 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[40]

	PIN DA[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 97.975 80.475 98.125 ;
			LAYER M2 ;
			RECT 80.295 97.975 80.475 98.125 ;
			LAYER M3 ;
			RECT 80.295 97.975 80.475 98.125 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[41]

	PIN DA[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 100.295 80.475 100.445 ;
			LAYER M2 ;
			RECT 80.295 100.295 80.475 100.445 ;
			LAYER M3 ;
			RECT 80.295 100.295 80.475 100.445 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[42]

	PIN DA[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 102.615 80.475 102.765 ;
			LAYER M1 ;
			RECT 80.295 102.615 80.475 102.765 ;
			LAYER M2 ;
			RECT 80.295 102.615 80.475 102.765 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[43]

	PIN DA[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 104.935 80.475 105.085 ;
			LAYER M2 ;
			RECT 80.295 104.935 80.475 105.085 ;
			LAYER M3 ;
			RECT 80.295 104.935 80.475 105.085 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[44]

	PIN DA[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 107.255 80.475 107.405 ;
			LAYER M1 ;
			RECT 80.295 107.255 80.475 107.405 ;
			LAYER M2 ;
			RECT 80.295 107.255 80.475 107.405 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[45]

	PIN DA[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 109.575 80.475 109.725 ;
			LAYER M1 ;
			RECT 80.295 109.575 80.475 109.725 ;
			LAYER M2 ;
			RECT 80.295 109.575 80.475 109.725 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[46]

	PIN DA[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 111.895 80.475 112.045 ;
			LAYER M2 ;
			RECT 80.295 111.895 80.475 112.045 ;
			LAYER M3 ;
			RECT 80.295 111.895 80.475 112.045 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[47]

	PIN DA[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 114.215 80.475 114.365 ;
			LAYER M2 ;
			RECT 80.295 114.215 80.475 114.365 ;
			LAYER M1 ;
			RECT 80.295 114.215 80.475 114.365 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[48]

	PIN DA[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 116.535 80.475 116.685 ;
			LAYER M3 ;
			RECT 80.295 116.535 80.475 116.685 ;
			LAYER M1 ;
			RECT 80.295 116.535 80.475 116.685 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[49]

	PIN DA[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 12.135 80.475 12.285 ;
			LAYER M1 ;
			RECT 80.295 12.135 80.475 12.285 ;
			LAYER M3 ;
			RECT 80.295 12.135 80.475 12.285 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[4]

	PIN DA[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 118.855 80.475 119.005 ;
			LAYER M2 ;
			RECT 80.295 118.855 80.475 119.005 ;
			LAYER M3 ;
			RECT 80.295 118.855 80.475 119.005 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[50]

	PIN DA[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 121.175 80.475 121.325 ;
			LAYER M1 ;
			RECT 80.295 121.175 80.475 121.325 ;
			LAYER M3 ;
			RECT 80.295 121.175 80.475 121.325 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[51]

	PIN DA[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 123.495 80.475 123.645 ;
			LAYER M1 ;
			RECT 80.295 123.495 80.475 123.645 ;
			LAYER M2 ;
			RECT 80.295 123.495 80.475 123.645 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[52]

	PIN DA[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 125.815 80.475 125.965 ;
			LAYER M2 ;
			RECT 80.295 125.815 80.475 125.965 ;
			LAYER M1 ;
			RECT 80.295 125.815 80.475 125.965 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[53]

	PIN DA[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 128.135 80.475 128.285 ;
			LAYER M1 ;
			RECT 80.295 128.135 80.475 128.285 ;
			LAYER M3 ;
			RECT 80.295 128.135 80.475 128.285 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[54]

	PIN DA[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 130.455 80.475 130.605 ;
			LAYER M2 ;
			RECT 80.295 130.455 80.475 130.605 ;
			LAYER M1 ;
			RECT 80.295 130.455 80.475 130.605 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[55]

	PIN DA[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 132.775 80.475 132.925 ;
			LAYER M1 ;
			RECT 80.295 132.775 80.475 132.925 ;
			LAYER M2 ;
			RECT 80.295 132.775 80.475 132.925 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[56]

	PIN DA[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 135.095 80.475 135.245 ;
			LAYER M2 ;
			RECT 80.295 135.095 80.475 135.245 ;
			LAYER M1 ;
			RECT 80.295 135.095 80.475 135.245 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[57]

	PIN DA[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 137.415 80.475 137.565 ;
			LAYER M3 ;
			RECT 80.295 137.415 80.475 137.565 ;
			LAYER M2 ;
			RECT 80.295 137.415 80.475 137.565 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[58]

	PIN DA[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 139.395 80.475 139.545 ;
			LAYER M3 ;
			RECT 80.295 139.395 80.475 139.545 ;
			LAYER M2 ;
			RECT 80.295 139.395 80.475 139.545 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[59]

	PIN DA[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 14.455 80.475 14.605 ;
			LAYER M2 ;
			RECT 80.295 14.455 80.475 14.605 ;
			LAYER M3 ;
			RECT 80.295 14.455 80.475 14.605 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[5]

	PIN DA[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 141.705 80.475 141.855 ;
			LAYER M1 ;
			RECT 80.295 141.705 80.475 141.855 ;
			LAYER M3 ;
			RECT 80.295 141.705 80.475 141.855 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[60]

	PIN DA[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 143.685 80.475 143.835 ;
			LAYER M1 ;
			RECT 80.295 143.685 80.475 143.835 ;
			LAYER M3 ;
			RECT 80.295 143.685 80.475 143.835 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[61]

	PIN DA[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 146.580 80.475 146.730 ;
			LAYER M1 ;
			RECT 80.295 146.580 80.475 146.730 ;
			LAYER M3 ;
			RECT 80.295 146.580 80.475 146.730 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[62]

	PIN DA[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 148.625 80.475 148.775 ;
			LAYER M2 ;
			RECT 80.295 148.625 80.475 148.775 ;
			LAYER M1 ;
			RECT 80.295 148.625 80.475 148.775 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[63]

	PIN DA[64]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 168.930 80.475 169.080 ;
			LAYER M3 ;
			RECT 80.295 168.930 80.475 169.080 ;
			LAYER M1 ;
			RECT 80.295 168.930 80.475 169.080 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[64]

	PIN DA[65]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 171.540 80.475 171.690 ;
			LAYER M1 ;
			RECT 80.295 171.540 80.475 171.690 ;
			LAYER M3 ;
			RECT 80.295 171.540 80.475 171.690 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[65]

	PIN DA[66]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 174.840 80.475 174.990 ;
			LAYER M2 ;
			RECT 80.295 174.840 80.475 174.990 ;
			LAYER M3 ;
			RECT 80.295 174.840 80.475 174.990 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[66]

	PIN DA[67]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 176.820 80.475 176.970 ;
			LAYER M3 ;
			RECT 80.295 176.820 80.475 176.970 ;
			LAYER M1 ;
			RECT 80.295 176.820 80.475 176.970 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[67]

	PIN DA[68]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 179.135 80.475 179.285 ;
			LAYER M2 ;
			RECT 80.295 179.135 80.475 179.285 ;
			LAYER M3 ;
			RECT 80.295 179.135 80.475 179.285 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[68]

	PIN DA[69]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 181.455 80.475 181.605 ;
			LAYER M1 ;
			RECT 80.295 181.455 80.475 181.605 ;
			LAYER M2 ;
			RECT 80.295 181.455 80.475 181.605 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[69]

	PIN DA[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 16.775 80.475 16.925 ;
			LAYER M1 ;
			RECT 80.295 16.775 80.475 16.925 ;
			LAYER M3 ;
			RECT 80.295 16.775 80.475 16.925 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[6]

	PIN DA[70]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 183.775 80.475 183.925 ;
			LAYER M1 ;
			RECT 80.295 183.775 80.475 183.925 ;
			LAYER M3 ;
			RECT 80.295 183.775 80.475 183.925 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[70]

	PIN DA[71]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 186.095 80.475 186.245 ;
			LAYER M2 ;
			RECT 80.295 186.095 80.475 186.245 ;
			LAYER M3 ;
			RECT 80.295 186.095 80.475 186.245 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[71]

	PIN DA[72]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 188.415 80.475 188.565 ;
			LAYER M2 ;
			RECT 80.295 188.415 80.475 188.565 ;
			LAYER M1 ;
			RECT 80.295 188.415 80.475 188.565 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[72]

	PIN DA[73]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 190.735 80.475 190.885 ;
			LAYER M2 ;
			RECT 80.295 190.735 80.475 190.885 ;
			LAYER M1 ;
			RECT 80.295 190.735 80.475 190.885 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[73]

	PIN DA[74]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 193.055 80.475 193.205 ;
			LAYER M3 ;
			RECT 80.295 193.055 80.475 193.205 ;
			LAYER M1 ;
			RECT 80.295 193.055 80.475 193.205 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[74]

	PIN DA[75]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 195.375 80.475 195.525 ;
			LAYER M3 ;
			RECT 80.295 195.375 80.475 195.525 ;
			LAYER M1 ;
			RECT 80.295 195.375 80.475 195.525 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[75]

	PIN DA[76]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 197.695 80.475 197.845 ;
			LAYER M1 ;
			RECT 80.295 197.695 80.475 197.845 ;
			LAYER M2 ;
			RECT 80.295 197.695 80.475 197.845 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[76]

	PIN DA[77]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 200.015 80.475 200.165 ;
			LAYER M2 ;
			RECT 80.295 200.015 80.475 200.165 ;
			LAYER M3 ;
			RECT 80.295 200.015 80.475 200.165 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[77]

	PIN DA[78]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 202.335 80.475 202.485 ;
			LAYER M1 ;
			RECT 80.295 202.335 80.475 202.485 ;
			LAYER M2 ;
			RECT 80.295 202.335 80.475 202.485 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[78]

	PIN DA[79]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 204.655 80.475 204.805 ;
			LAYER M2 ;
			RECT 80.295 204.655 80.475 204.805 ;
			LAYER M3 ;
			RECT 80.295 204.655 80.475 204.805 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[79]

	PIN DA[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 19.095 80.475 19.245 ;
			LAYER M2 ;
			RECT 80.295 19.095 80.475 19.245 ;
			LAYER M1 ;
			RECT 80.295 19.095 80.475 19.245 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[7]

	PIN DA[80]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 206.975 80.475 207.125 ;
			LAYER M2 ;
			RECT 80.295 206.975 80.475 207.125 ;
			LAYER M3 ;
			RECT 80.295 206.975 80.475 207.125 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[80]

	PIN DA[81]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 209.295 80.475 209.445 ;
			LAYER M3 ;
			RECT 80.295 209.295 80.475 209.445 ;
			LAYER M1 ;
			RECT 80.295 209.295 80.475 209.445 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[81]

	PIN DA[82]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 211.615 80.475 211.765 ;
			LAYER M1 ;
			RECT 80.295 211.615 80.475 211.765 ;
			LAYER M3 ;
			RECT 80.295 211.615 80.475 211.765 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[82]

	PIN DA[83]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 213.935 80.475 214.085 ;
			LAYER M1 ;
			RECT 80.295 213.935 80.475 214.085 ;
			LAYER M2 ;
			RECT 80.295 213.935 80.475 214.085 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[83]

	PIN DA[84]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 216.255 80.475 216.405 ;
			LAYER M2 ;
			RECT 80.295 216.255 80.475 216.405 ;
			LAYER M3 ;
			RECT 80.295 216.255 80.475 216.405 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[84]

	PIN DA[85]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 218.575 80.475 218.725 ;
			LAYER M3 ;
			RECT 80.295 218.575 80.475 218.725 ;
			LAYER M2 ;
			RECT 80.295 218.575 80.475 218.725 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[85]

	PIN DA[86]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 220.895 80.475 221.045 ;
			LAYER M3 ;
			RECT 80.295 220.895 80.475 221.045 ;
			LAYER M1 ;
			RECT 80.295 220.895 80.475 221.045 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[86]

	PIN DA[87]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 223.215 80.475 223.365 ;
			LAYER M2 ;
			RECT 80.295 223.215 80.475 223.365 ;
			LAYER M1 ;
			RECT 80.295 223.215 80.475 223.365 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[87]

	PIN DA[88]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 225.535 80.475 225.685 ;
			LAYER M3 ;
			RECT 80.295 225.535 80.475 225.685 ;
			LAYER M2 ;
			RECT 80.295 225.535 80.475 225.685 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[88]

	PIN DA[89]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 227.855 80.475 228.005 ;
			LAYER M1 ;
			RECT 80.295 227.855 80.475 228.005 ;
			LAYER M3 ;
			RECT 80.295 227.855 80.475 228.005 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[89]

	PIN DA[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 21.415 80.475 21.565 ;
			LAYER M3 ;
			RECT 80.295 21.415 80.475 21.565 ;
			LAYER M2 ;
			RECT 80.295 21.415 80.475 21.565 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[8]

	PIN DA[90]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 230.175 80.475 230.325 ;
			LAYER M2 ;
			RECT 80.295 230.175 80.475 230.325 ;
			LAYER M1 ;
			RECT 80.295 230.175 80.475 230.325 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[90]

	PIN DA[91]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 232.495 80.475 232.645 ;
			LAYER M1 ;
			RECT 80.295 232.495 80.475 232.645 ;
			LAYER M2 ;
			RECT 80.295 232.495 80.475 232.645 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[91]

	PIN DA[92]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 234.815 80.475 234.965 ;
			LAYER M2 ;
			RECT 80.295 234.815 80.475 234.965 ;
			LAYER M3 ;
			RECT 80.295 234.815 80.475 234.965 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[92]

	PIN DA[93]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 237.135 80.475 237.285 ;
			LAYER M1 ;
			RECT 80.295 237.135 80.475 237.285 ;
			LAYER M3 ;
			RECT 80.295 237.135 80.475 237.285 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[93]

	PIN DA[94]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 239.455 80.475 239.605 ;
			LAYER M2 ;
			RECT 80.295 239.455 80.475 239.605 ;
			LAYER M3 ;
			RECT 80.295 239.455 80.475 239.605 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[94]

	PIN DA[95]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 241.775 80.475 241.925 ;
			LAYER M1 ;
			RECT 80.295 241.775 80.475 241.925 ;
			LAYER M2 ;
			RECT 80.295 241.775 80.475 241.925 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[95]

	PIN DA[96]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 244.095 80.475 244.245 ;
			LAYER M1 ;
			RECT 80.295 244.095 80.475 244.245 ;
			LAYER M2 ;
			RECT 80.295 244.095 80.475 244.245 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[96]

	PIN DA[97]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 246.415 80.475 246.565 ;
			LAYER M1 ;
			RECT 80.295 246.415 80.475 246.565 ;
			LAYER M3 ;
			RECT 80.295 246.415 80.475 246.565 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[97]

	PIN DA[98]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 248.735 80.475 248.885 ;
			LAYER M3 ;
			RECT 80.295 248.735 80.475 248.885 ;
			LAYER M1 ;
			RECT 80.295 248.735 80.475 248.885 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[98]

	PIN DA[99]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 251.055 80.475 251.205 ;
			LAYER M2 ;
			RECT 80.295 251.055 80.475 251.205 ;
			LAYER M1 ;
			RECT 80.295 251.055 80.475 251.205 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[99]

	PIN DA[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 23.735 80.475 23.885 ;
			LAYER M2 ;
			RECT 80.295 23.735 80.475 23.885 ;
			LAYER M3 ;
			RECT 80.295 23.735 80.475 23.885 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[9]

	PIN DB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 3.185 80.475 3.335 ;
			LAYER M1 ;
			RECT 80.295 3.185 80.475 3.335 ;
			LAYER M3 ;
			RECT 80.295 3.185 80.475 3.335 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[0]

	PIN DB[100]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 253.705 80.475 253.855 ;
			LAYER M2 ;
			RECT 80.295 253.705 80.475 253.855 ;
			LAYER M1 ;
			RECT 80.295 253.705 80.475 253.855 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[100]

	PIN DB[101]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 256.025 80.475 256.175 ;
			LAYER M2 ;
			RECT 80.295 256.025 80.475 256.175 ;
			LAYER M3 ;
			RECT 80.295 256.025 80.475 256.175 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[101]

	PIN DB[102]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 258.345 80.475 258.495 ;
			LAYER M3 ;
			RECT 80.295 258.345 80.475 258.495 ;
			LAYER M2 ;
			RECT 80.295 258.345 80.475 258.495 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[102]

	PIN DB[103]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 260.665 80.475 260.815 ;
			LAYER M2 ;
			RECT 80.295 260.665 80.475 260.815 ;
			LAYER M1 ;
			RECT 80.295 260.665 80.475 260.815 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[103]

	PIN DB[104]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 262.985 80.475 263.135 ;
			LAYER M3 ;
			RECT 80.295 262.985 80.475 263.135 ;
			LAYER M1 ;
			RECT 80.295 262.985 80.475 263.135 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[104]

	PIN DB[105]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 265.305 80.475 265.455 ;
			LAYER M3 ;
			RECT 80.295 265.305 80.475 265.455 ;
			LAYER M2 ;
			RECT 80.295 265.305 80.475 265.455 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[105]

	PIN DB[106]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 267.625 80.475 267.775 ;
			LAYER M2 ;
			RECT 80.295 267.625 80.475 267.775 ;
			LAYER M1 ;
			RECT 80.295 267.625 80.475 267.775 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[106]

	PIN DB[107]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 269.945 80.475 270.095 ;
			LAYER M1 ;
			RECT 80.295 269.945 80.475 270.095 ;
			LAYER M2 ;
			RECT 80.295 269.945 80.475 270.095 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[107]

	PIN DB[108]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 272.265 80.475 272.415 ;
			LAYER M2 ;
			RECT 80.295 272.265 80.475 272.415 ;
			LAYER M1 ;
			RECT 80.295 272.265 80.475 272.415 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[108]

	PIN DB[109]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 274.585 80.475 274.735 ;
			LAYER M2 ;
			RECT 80.295 274.585 80.475 274.735 ;
			LAYER M3 ;
			RECT 80.295 274.585 80.475 274.735 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[109]

	PIN DB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 26.385 80.475 26.535 ;
			LAYER M3 ;
			RECT 80.295 26.385 80.475 26.535 ;
			LAYER M2 ;
			RECT 80.295 26.385 80.475 26.535 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[10]

	PIN DB[110]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 276.905 80.475 277.055 ;
			LAYER M2 ;
			RECT 80.295 276.905 80.475 277.055 ;
			LAYER M1 ;
			RECT 80.295 276.905 80.475 277.055 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[110]

	PIN DB[111]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 279.225 80.475 279.375 ;
			LAYER M2 ;
			RECT 80.295 279.225 80.475 279.375 ;
			LAYER M1 ;
			RECT 80.295 279.225 80.475 279.375 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[111]

	PIN DB[112]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 281.545 80.475 281.695 ;
			LAYER M3 ;
			RECT 80.295 281.545 80.475 281.695 ;
			LAYER M1 ;
			RECT 80.295 281.545 80.475 281.695 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[112]

	PIN DB[113]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 283.865 80.475 284.015 ;
			LAYER M3 ;
			RECT 80.295 283.865 80.475 284.015 ;
			LAYER M2 ;
			RECT 80.295 283.865 80.475 284.015 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[113]

	PIN DB[114]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 286.185 80.475 286.335 ;
			LAYER M3 ;
			RECT 80.295 286.185 80.475 286.335 ;
			LAYER M2 ;
			RECT 80.295 286.185 80.475 286.335 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[114]

	PIN DB[115]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 288.505 80.475 288.655 ;
			LAYER M1 ;
			RECT 80.295 288.505 80.475 288.655 ;
			LAYER M3 ;
			RECT 80.295 288.505 80.475 288.655 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[115]

	PIN DB[116]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 290.825 80.475 290.975 ;
			LAYER M2 ;
			RECT 80.295 290.825 80.475 290.975 ;
			LAYER M1 ;
			RECT 80.295 290.825 80.475 290.975 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[116]

	PIN DB[117]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 293.145 80.475 293.295 ;
			LAYER M2 ;
			RECT 80.295 293.145 80.475 293.295 ;
			LAYER M1 ;
			RECT 80.295 293.145 80.475 293.295 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[117]

	PIN DB[118]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 295.465 80.475 295.615 ;
			LAYER M3 ;
			RECT 80.295 295.465 80.475 295.615 ;
			LAYER M1 ;
			RECT 80.295 295.465 80.475 295.615 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[118]

	PIN DB[119]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 297.785 80.475 297.935 ;
			LAYER M1 ;
			RECT 80.295 297.785 80.475 297.935 ;
			LAYER M2 ;
			RECT 80.295 297.785 80.475 297.935 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[119]

	PIN DB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 28.705 80.475 28.855 ;
			LAYER M3 ;
			RECT 80.295 28.705 80.475 28.855 ;
			LAYER M2 ;
			RECT 80.295 28.705 80.475 28.855 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[11]

	PIN DB[120]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 300.105 80.475 300.255 ;
			LAYER M3 ;
			RECT 80.295 300.105 80.475 300.255 ;
			LAYER M1 ;
			RECT 80.295 300.105 80.475 300.255 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[120]

	PIN DB[121]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 302.425 80.475 302.575 ;
			LAYER M1 ;
			RECT 80.295 302.425 80.475 302.575 ;
			LAYER M3 ;
			RECT 80.295 302.425 80.475 302.575 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[121]

	PIN DB[122]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 304.745 80.475 304.895 ;
			LAYER M2 ;
			RECT 80.295 304.745 80.475 304.895 ;
			LAYER M1 ;
			RECT 80.295 304.745 80.475 304.895 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[122]

	PIN DB[123]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 307.065 80.475 307.215 ;
			LAYER M1 ;
			RECT 80.295 307.065 80.475 307.215 ;
			LAYER M3 ;
			RECT 80.295 307.065 80.475 307.215 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[123]

	PIN DB[124]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 309.385 80.475 309.535 ;
			LAYER M1 ;
			RECT 80.295 309.385 80.475 309.535 ;
			LAYER M3 ;
			RECT 80.295 309.385 80.475 309.535 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[124]

	PIN DB[125]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 311.705 80.475 311.855 ;
			LAYER M2 ;
			RECT 80.295 311.705 80.475 311.855 ;
			LAYER M1 ;
			RECT 80.295 311.705 80.475 311.855 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[125]

	PIN DB[126]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 314.025 80.475 314.175 ;
			LAYER M2 ;
			RECT 80.295 314.025 80.475 314.175 ;
			LAYER M1 ;
			RECT 80.295 314.025 80.475 314.175 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[126]

	PIN DB[127]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 316.345 80.475 316.495 ;
			LAYER M2 ;
			RECT 80.295 316.345 80.475 316.495 ;
			LAYER M3 ;
			RECT 80.295 316.345 80.475 316.495 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[127]

	PIN DB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 31.025 80.475 31.175 ;
			LAYER M1 ;
			RECT 80.295 31.025 80.475 31.175 ;
			LAYER M3 ;
			RECT 80.295 31.025 80.475 31.175 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[12]

	PIN DB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 33.345 80.475 33.495 ;
			LAYER M1 ;
			RECT 80.295 33.345 80.475 33.495 ;
			LAYER M3 ;
			RECT 80.295 33.345 80.475 33.495 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[13]

	PIN DB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 35.665 80.475 35.815 ;
			LAYER M1 ;
			RECT 80.295 35.665 80.475 35.815 ;
			LAYER M2 ;
			RECT 80.295 35.665 80.475 35.815 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[14]

	PIN DB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 37.985 80.475 38.135 ;
			LAYER M2 ;
			RECT 80.295 37.985 80.475 38.135 ;
			LAYER M1 ;
			RECT 80.295 37.985 80.475 38.135 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[15]

	PIN DB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 40.305 80.475 40.455 ;
			LAYER M2 ;
			RECT 80.295 40.305 80.475 40.455 ;
			LAYER M1 ;
			RECT 80.295 40.305 80.475 40.455 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[16]

	PIN DB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 42.625 80.475 42.775 ;
			LAYER M2 ;
			RECT 80.295 42.625 80.475 42.775 ;
			LAYER M1 ;
			RECT 80.295 42.625 80.475 42.775 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[17]

	PIN DB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 44.945 80.475 45.095 ;
			LAYER M1 ;
			RECT 80.295 44.945 80.475 45.095 ;
			LAYER M3 ;
			RECT 80.295 44.945 80.475 45.095 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[18]

	PIN DB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 47.265 80.475 47.415 ;
			LAYER M2 ;
			RECT 80.295 47.265 80.475 47.415 ;
			LAYER M1 ;
			RECT 80.295 47.265 80.475 47.415 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[19]

	PIN DB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 5.505 80.475 5.655 ;
			LAYER M3 ;
			RECT 80.295 5.505 80.475 5.655 ;
			LAYER M1 ;
			RECT 80.295 5.505 80.475 5.655 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[1]

	PIN DB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 49.585 80.475 49.735 ;
			LAYER M3 ;
			RECT 80.295 49.585 80.475 49.735 ;
			LAYER M2 ;
			RECT 80.295 49.585 80.475 49.735 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[20]

	PIN DB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 51.905 80.475 52.055 ;
			LAYER M1 ;
			RECT 80.295 51.905 80.475 52.055 ;
			LAYER M2 ;
			RECT 80.295 51.905 80.475 52.055 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[21]

	PIN DB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 54.225 80.475 54.375 ;
			LAYER M2 ;
			RECT 80.295 54.225 80.475 54.375 ;
			LAYER M1 ;
			RECT 80.295 54.225 80.475 54.375 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[22]

	PIN DB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 56.545 80.475 56.695 ;
			LAYER M2 ;
			RECT 80.295 56.545 80.475 56.695 ;
			LAYER M1 ;
			RECT 80.295 56.545 80.475 56.695 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[23]

	PIN DB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 58.865 80.475 59.015 ;
			LAYER M2 ;
			RECT 80.295 58.865 80.475 59.015 ;
			LAYER M3 ;
			RECT 80.295 58.865 80.475 59.015 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[24]

	PIN DB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 61.185 80.475 61.335 ;
			LAYER M1 ;
			RECT 80.295 61.185 80.475 61.335 ;
			LAYER M3 ;
			RECT 80.295 61.185 80.475 61.335 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[25]

	PIN DB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 63.505 80.475 63.655 ;
			LAYER M1 ;
			RECT 80.295 63.505 80.475 63.655 ;
			LAYER M2 ;
			RECT 80.295 63.505 80.475 63.655 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[26]

	PIN DB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 65.825 80.475 65.975 ;
			LAYER M3 ;
			RECT 80.295 65.825 80.475 65.975 ;
			LAYER M1 ;
			RECT 80.295 65.825 80.475 65.975 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[27]

	PIN DB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 68.145 80.475 68.295 ;
			LAYER M2 ;
			RECT 80.295 68.145 80.475 68.295 ;
			LAYER M1 ;
			RECT 80.295 68.145 80.475 68.295 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[28]

	PIN DB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 70.465 80.475 70.615 ;
			LAYER M1 ;
			RECT 80.295 70.465 80.475 70.615 ;
			LAYER M3 ;
			RECT 80.295 70.465 80.475 70.615 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[29]

	PIN DB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 7.825 80.475 7.975 ;
			LAYER M2 ;
			RECT 80.295 7.825 80.475 7.975 ;
			LAYER M1 ;
			RECT 80.295 7.825 80.475 7.975 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[2]

	PIN DB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 72.785 80.475 72.935 ;
			LAYER M1 ;
			RECT 80.295 72.785 80.475 72.935 ;
			LAYER M3 ;
			RECT 80.295 72.785 80.475 72.935 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[30]

	PIN DB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 75.105 80.475 75.255 ;
			LAYER M1 ;
			RECT 80.295 75.105 80.475 75.255 ;
			LAYER M3 ;
			RECT 80.295 75.105 80.475 75.255 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[31]

	PIN DB[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 77.425 80.475 77.575 ;
			LAYER M3 ;
			RECT 80.295 77.425 80.475 77.575 ;
			LAYER M1 ;
			RECT 80.295 77.425 80.475 77.575 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[32]

	PIN DB[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 79.745 80.475 79.895 ;
			LAYER M2 ;
			RECT 80.295 79.745 80.475 79.895 ;
			LAYER M3 ;
			RECT 80.295 79.745 80.475 79.895 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[33]

	PIN DB[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 82.065 80.475 82.215 ;
			LAYER M1 ;
			RECT 80.295 82.065 80.475 82.215 ;
			LAYER M2 ;
			RECT 80.295 82.065 80.475 82.215 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[34]

	PIN DB[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 84.385 80.475 84.535 ;
			LAYER M3 ;
			RECT 80.295 84.385 80.475 84.535 ;
			LAYER M1 ;
			RECT 80.295 84.385 80.475 84.535 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[35]

	PIN DB[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 86.705 80.475 86.855 ;
			LAYER M1 ;
			RECT 80.295 86.705 80.475 86.855 ;
			LAYER M3 ;
			RECT 80.295 86.705 80.475 86.855 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[36]

	PIN DB[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 89.025 80.475 89.175 ;
			LAYER M1 ;
			RECT 80.295 89.025 80.475 89.175 ;
			LAYER M3 ;
			RECT 80.295 89.025 80.475 89.175 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[37]

	PIN DB[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 91.345 80.475 91.495 ;
			LAYER M3 ;
			RECT 80.295 91.345 80.475 91.495 ;
			LAYER M2 ;
			RECT 80.295 91.345 80.475 91.495 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[38]

	PIN DB[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 93.665 80.475 93.815 ;
			LAYER M1 ;
			RECT 80.295 93.665 80.475 93.815 ;
			LAYER M3 ;
			RECT 80.295 93.665 80.475 93.815 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[39]

	PIN DB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 10.145 80.475 10.295 ;
			LAYER M2 ;
			RECT 80.295 10.145 80.475 10.295 ;
			LAYER M1 ;
			RECT 80.295 10.145 80.475 10.295 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[3]

	PIN DB[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 95.985 80.475 96.135 ;
			LAYER M2 ;
			RECT 80.295 95.985 80.475 96.135 ;
			LAYER M1 ;
			RECT 80.295 95.985 80.475 96.135 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[40]

	PIN DB[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 98.305 80.475 98.455 ;
			LAYER M2 ;
			RECT 80.295 98.305 80.475 98.455 ;
			LAYER M1 ;
			RECT 80.295 98.305 80.475 98.455 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[41]

	PIN DB[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 100.625 80.475 100.775 ;
			LAYER M1 ;
			RECT 80.295 100.625 80.475 100.775 ;
			LAYER M3 ;
			RECT 80.295 100.625 80.475 100.775 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[42]

	PIN DB[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 102.945 80.475 103.095 ;
			LAYER M1 ;
			RECT 80.295 102.945 80.475 103.095 ;
			LAYER M2 ;
			RECT 80.295 102.945 80.475 103.095 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[43]

	PIN DB[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 105.265 80.475 105.415 ;
			LAYER M2 ;
			RECT 80.295 105.265 80.475 105.415 ;
			LAYER M1 ;
			RECT 80.295 105.265 80.475 105.415 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[44]

	PIN DB[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 107.585 80.475 107.735 ;
			LAYER M1 ;
			RECT 80.295 107.585 80.475 107.735 ;
			LAYER M2 ;
			RECT 80.295 107.585 80.475 107.735 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[45]

	PIN DB[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 109.905 80.475 110.055 ;
			LAYER M2 ;
			RECT 80.295 109.905 80.475 110.055 ;
			LAYER M1 ;
			RECT 80.295 109.905 80.475 110.055 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[46]

	PIN DB[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 112.225 80.475 112.375 ;
			LAYER M3 ;
			RECT 80.295 112.225 80.475 112.375 ;
			LAYER M1 ;
			RECT 80.295 112.225 80.475 112.375 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[47]

	PIN DB[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 114.545 80.475 114.695 ;
			LAYER M1 ;
			RECT 80.295 114.545 80.475 114.695 ;
			LAYER M3 ;
			RECT 80.295 114.545 80.475 114.695 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[48]

	PIN DB[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 116.865 80.475 117.015 ;
			LAYER M1 ;
			RECT 80.295 116.865 80.475 117.015 ;
			LAYER M3 ;
			RECT 80.295 116.865 80.475 117.015 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[49]

	PIN DB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 12.465 80.475 12.615 ;
			LAYER M3 ;
			RECT 80.295 12.465 80.475 12.615 ;
			LAYER M2 ;
			RECT 80.295 12.465 80.475 12.615 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[4]

	PIN DB[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 119.185 80.475 119.335 ;
			LAYER M3 ;
			RECT 80.295 119.185 80.475 119.335 ;
			LAYER M1 ;
			RECT 80.295 119.185 80.475 119.335 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[50]

	PIN DB[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 121.505 80.475 121.655 ;
			LAYER M2 ;
			RECT 80.295 121.505 80.475 121.655 ;
			LAYER M1 ;
			RECT 80.295 121.505 80.475 121.655 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[51]

	PIN DB[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 123.825 80.475 123.975 ;
			LAYER M1 ;
			RECT 80.295 123.825 80.475 123.975 ;
			LAYER M3 ;
			RECT 80.295 123.825 80.475 123.975 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[52]

	PIN DB[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 126.145 80.475 126.295 ;
			LAYER M3 ;
			RECT 80.295 126.145 80.475 126.295 ;
			LAYER M1 ;
			RECT 80.295 126.145 80.475 126.295 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[53]

	PIN DB[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 128.465 80.475 128.615 ;
			LAYER M1 ;
			RECT 80.295 128.465 80.475 128.615 ;
			LAYER M3 ;
			RECT 80.295 128.465 80.475 128.615 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[54]

	PIN DB[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 130.785 80.475 130.935 ;
			LAYER M2 ;
			RECT 80.295 130.785 80.475 130.935 ;
			LAYER M1 ;
			RECT 80.295 130.785 80.475 130.935 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[55]

	PIN DB[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 133.105 80.475 133.255 ;
			LAYER M2 ;
			RECT 80.295 133.105 80.475 133.255 ;
			LAYER M1 ;
			RECT 80.295 133.105 80.475 133.255 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[56]

	PIN DB[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 135.425 80.475 135.575 ;
			LAYER M1 ;
			RECT 80.295 135.425 80.475 135.575 ;
			LAYER M3 ;
			RECT 80.295 135.425 80.475 135.575 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[57]

	PIN DB[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 137.745 80.475 137.895 ;
			LAYER M2 ;
			RECT 80.295 137.745 80.475 137.895 ;
			LAYER M3 ;
			RECT 80.295 137.745 80.475 137.895 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[58]

	PIN DB[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 140.055 80.475 140.205 ;
			LAYER M3 ;
			RECT 80.295 140.055 80.475 140.205 ;
			LAYER M1 ;
			RECT 80.295 140.055 80.475 140.205 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[59]

	PIN DB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 14.785 80.475 14.935 ;
			LAYER M3 ;
			RECT 80.295 14.785 80.475 14.935 ;
			LAYER M2 ;
			RECT 80.295 14.785 80.475 14.935 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[5]

	PIN DB[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 142.035 80.475 142.185 ;
			LAYER M2 ;
			RECT 80.295 142.035 80.475 142.185 ;
			LAYER M1 ;
			RECT 80.295 142.035 80.475 142.185 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[60]

	PIN DB[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 144.930 80.475 145.080 ;
			LAYER M2 ;
			RECT 80.295 144.930 80.475 145.080 ;
			LAYER M3 ;
			RECT 80.295 144.930 80.475 145.080 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[61]

	PIN DB[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 146.910 80.475 147.060 ;
			LAYER M3 ;
			RECT 80.295 146.910 80.475 147.060 ;
			LAYER M1 ;
			RECT 80.295 146.910 80.475 147.060 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[62]

	PIN DB[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 148.955 80.475 149.105 ;
			LAYER M2 ;
			RECT 80.295 148.955 80.475 149.105 ;
			LAYER M1 ;
			RECT 80.295 148.955 80.475 149.105 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[63]

	PIN DB[64]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 169.890 80.475 170.040 ;
			LAYER M1 ;
			RECT 80.295 169.890 80.475 170.040 ;
			LAYER M3 ;
			RECT 80.295 169.890 80.475 170.040 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[64]

	PIN DB[65]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 172.200 80.475 172.350 ;
			LAYER M1 ;
			RECT 80.295 172.200 80.475 172.350 ;
			LAYER M3 ;
			RECT 80.295 172.200 80.475 172.350 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[65]

	PIN DB[66]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 175.170 80.475 175.320 ;
			LAYER M2 ;
			RECT 80.295 175.170 80.475 175.320 ;
			LAYER M3 ;
			RECT 80.295 175.170 80.475 175.320 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[66]

	PIN DB[67]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 177.480 80.475 177.630 ;
			LAYER M2 ;
			RECT 80.295 177.480 80.475 177.630 ;
			LAYER M1 ;
			RECT 80.295 177.480 80.475 177.630 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[67]

	PIN DB[68]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 179.465 80.475 179.615 ;
			LAYER M3 ;
			RECT 80.295 179.465 80.475 179.615 ;
			LAYER M1 ;
			RECT 80.295 179.465 80.475 179.615 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[68]

	PIN DB[69]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 181.785 80.475 181.935 ;
			LAYER M2 ;
			RECT 80.295 181.785 80.475 181.935 ;
			LAYER M1 ;
			RECT 80.295 181.785 80.475 181.935 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[69]

	PIN DB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 17.105 80.475 17.255 ;
			LAYER M2 ;
			RECT 80.295 17.105 80.475 17.255 ;
			LAYER M3 ;
			RECT 80.295 17.105 80.475 17.255 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[6]

	PIN DB[70]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 184.105 80.475 184.255 ;
			LAYER M1 ;
			RECT 80.295 184.105 80.475 184.255 ;
			LAYER M2 ;
			RECT 80.295 184.105 80.475 184.255 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[70]

	PIN DB[71]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 186.425 80.475 186.575 ;
			LAYER M2 ;
			RECT 80.295 186.425 80.475 186.575 ;
			LAYER M3 ;
			RECT 80.295 186.425 80.475 186.575 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[71]

	PIN DB[72]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 188.745 80.475 188.895 ;
			LAYER M3 ;
			RECT 80.295 188.745 80.475 188.895 ;
			LAYER M2 ;
			RECT 80.295 188.745 80.475 188.895 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[72]

	PIN DB[73]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 191.065 80.475 191.215 ;
			LAYER M1 ;
			RECT 80.295 191.065 80.475 191.215 ;
			LAYER M2 ;
			RECT 80.295 191.065 80.475 191.215 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[73]

	PIN DB[74]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 193.385 80.475 193.535 ;
			LAYER M1 ;
			RECT 80.295 193.385 80.475 193.535 ;
			LAYER M2 ;
			RECT 80.295 193.385 80.475 193.535 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[74]

	PIN DB[75]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 195.705 80.475 195.855 ;
			LAYER M3 ;
			RECT 80.295 195.705 80.475 195.855 ;
			LAYER M2 ;
			RECT 80.295 195.705 80.475 195.855 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[75]

	PIN DB[76]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 198.025 80.475 198.175 ;
			LAYER M2 ;
			RECT 80.295 198.025 80.475 198.175 ;
			LAYER M1 ;
			RECT 80.295 198.025 80.475 198.175 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[76]

	PIN DB[77]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 200.345 80.475 200.495 ;
			LAYER M1 ;
			RECT 80.295 200.345 80.475 200.495 ;
			LAYER M2 ;
			RECT 80.295 200.345 80.475 200.495 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[77]

	PIN DB[78]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 202.665 80.475 202.815 ;
			LAYER M1 ;
			RECT 80.295 202.665 80.475 202.815 ;
			LAYER M3 ;
			RECT 80.295 202.665 80.475 202.815 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[78]

	PIN DB[79]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 204.985 80.475 205.135 ;
			LAYER M2 ;
			RECT 80.295 204.985 80.475 205.135 ;
			LAYER M1 ;
			RECT 80.295 204.985 80.475 205.135 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[79]

	PIN DB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 19.425 80.475 19.575 ;
			LAYER M3 ;
			RECT 80.295 19.425 80.475 19.575 ;
			LAYER M1 ;
			RECT 80.295 19.425 80.475 19.575 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[7]

	PIN DB[80]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 207.305 80.475 207.455 ;
			LAYER M2 ;
			RECT 80.295 207.305 80.475 207.455 ;
			LAYER M3 ;
			RECT 80.295 207.305 80.475 207.455 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[80]

	PIN DB[81]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 209.625 80.475 209.775 ;
			LAYER M2 ;
			RECT 80.295 209.625 80.475 209.775 ;
			LAYER M1 ;
			RECT 80.295 209.625 80.475 209.775 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[81]

	PIN DB[82]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 211.945 80.475 212.095 ;
			LAYER M2 ;
			RECT 80.295 211.945 80.475 212.095 ;
			LAYER M1 ;
			RECT 80.295 211.945 80.475 212.095 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[82]

	PIN DB[83]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 214.265 80.475 214.415 ;
			LAYER M1 ;
			RECT 80.295 214.265 80.475 214.415 ;
			LAYER M2 ;
			RECT 80.295 214.265 80.475 214.415 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[83]

	PIN DB[84]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 216.585 80.475 216.735 ;
			LAYER M2 ;
			RECT 80.295 216.585 80.475 216.735 ;
			LAYER M3 ;
			RECT 80.295 216.585 80.475 216.735 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[84]

	PIN DB[85]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 218.905 80.475 219.055 ;
			LAYER M1 ;
			RECT 80.295 218.905 80.475 219.055 ;
			LAYER M3 ;
			RECT 80.295 218.905 80.475 219.055 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[85]

	PIN DB[86]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 221.225 80.475 221.375 ;
			LAYER M1 ;
			RECT 80.295 221.225 80.475 221.375 ;
			LAYER M3 ;
			RECT 80.295 221.225 80.475 221.375 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[86]

	PIN DB[87]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 223.545 80.475 223.695 ;
			LAYER M3 ;
			RECT 80.295 223.545 80.475 223.695 ;
			LAYER M1 ;
			RECT 80.295 223.545 80.475 223.695 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[87]

	PIN DB[88]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 225.865 80.475 226.015 ;
			LAYER M2 ;
			RECT 80.295 225.865 80.475 226.015 ;
			LAYER M3 ;
			RECT 80.295 225.865 80.475 226.015 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[88]

	PIN DB[89]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 228.185 80.475 228.335 ;
			LAYER M2 ;
			RECT 80.295 228.185 80.475 228.335 ;
			LAYER M3 ;
			RECT 80.295 228.185 80.475 228.335 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[89]

	PIN DB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 21.745 80.475 21.895 ;
			LAYER M2 ;
			RECT 80.295 21.745 80.475 21.895 ;
			LAYER M1 ;
			RECT 80.295 21.745 80.475 21.895 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[8]

	PIN DB[90]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 230.505 80.475 230.655 ;
			LAYER M2 ;
			RECT 80.295 230.505 80.475 230.655 ;
			LAYER M3 ;
			RECT 80.295 230.505 80.475 230.655 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[90]

	PIN DB[91]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 232.825 80.475 232.975 ;
			LAYER M2 ;
			RECT 80.295 232.825 80.475 232.975 ;
			LAYER M3 ;
			RECT 80.295 232.825 80.475 232.975 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[91]

	PIN DB[92]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 235.145 80.475 235.295 ;
			LAYER M2 ;
			RECT 80.295 235.145 80.475 235.295 ;
			LAYER M1 ;
			RECT 80.295 235.145 80.475 235.295 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[92]

	PIN DB[93]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 237.465 80.475 237.615 ;
			LAYER M3 ;
			RECT 80.295 237.465 80.475 237.615 ;
			LAYER M1 ;
			RECT 80.295 237.465 80.475 237.615 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[93]

	PIN DB[94]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 239.785 80.475 239.935 ;
			LAYER M3 ;
			RECT 80.295 239.785 80.475 239.935 ;
			LAYER M2 ;
			RECT 80.295 239.785 80.475 239.935 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[94]

	PIN DB[95]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 242.105 80.475 242.255 ;
			LAYER M2 ;
			RECT 80.295 242.105 80.475 242.255 ;
			LAYER M1 ;
			RECT 80.295 242.105 80.475 242.255 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[95]

	PIN DB[96]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 244.425 80.475 244.575 ;
			LAYER M1 ;
			RECT 80.295 244.425 80.475 244.575 ;
			LAYER M2 ;
			RECT 80.295 244.425 80.475 244.575 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[96]

	PIN DB[97]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 246.745 80.475 246.895 ;
			LAYER M3 ;
			RECT 80.295 246.745 80.475 246.895 ;
			LAYER M1 ;
			RECT 80.295 246.745 80.475 246.895 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[97]

	PIN DB[98]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 249.065 80.475 249.215 ;
			LAYER M1 ;
			RECT 80.295 249.065 80.475 249.215 ;
			LAYER M3 ;
			RECT 80.295 249.065 80.475 249.215 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[98]

	PIN DB[99]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 251.385 80.475 251.535 ;
			LAYER M1 ;
			RECT 80.295 251.385 80.475 251.535 ;
			LAYER M2 ;
			RECT 80.295 251.385 80.475 251.535 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[99]

	PIN DB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 24.065 80.475 24.215 ;
			LAYER M1 ;
			RECT 80.295 24.065 80.475 24.215 ;
			LAYER M3 ;
			RECT 80.295 24.065 80.475 24.215 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[9]

	PIN PTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 163.980 80.475 164.130 ;
			LAYER M2 ;
			RECT 80.295 163.980 80.475 164.130 ;
			LAYER M3 ;
			RECT 80.295 163.980 80.475 164.130 ;
		END
		ANTENNAGATEAREA 0.015900 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.219900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.012600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.408800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.015900 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483500 LAYER M2 ;
		ANTENNAMAXAREACAR 31.421400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.817600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.015900 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121200 LAYER M3 ;
		ANTENNAMAXAREACAR 33.119500 LAYER M3 ;
	END PTSEL[0]

	PIN PTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 164.310 80.475 164.460 ;
			LAYER M3 ;
			RECT 80.295 164.310 80.475 164.460 ;
			LAYER M1 ;
			RECT 80.295 164.310 80.475 164.460 ;
		END
		ANTENNAGATEAREA 0.015900 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.219900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.012600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.408800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.015900 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483500 LAYER M2 ;
		ANTENNAMAXAREACAR 31.421400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.817600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.015900 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121200 LAYER M3 ;
		ANTENNAMAXAREACAR 33.119500 LAYER M3 ;
	END PTSEL[1]

	PIN QA[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 1.860 80.475 2.010 ;
			LAYER M3 ;
			RECT 80.295 1.860 80.475 2.010 ;
			LAYER M1 ;
			RECT 80.295 1.860 80.475 2.010 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[0]

	PIN QA[100]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 252.380 80.475 252.530 ;
			LAYER M1 ;
			RECT 80.295 252.380 80.475 252.530 ;
			LAYER M2 ;
			RECT 80.295 252.380 80.475 252.530 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[100]

	PIN QA[101]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 254.700 80.475 254.850 ;
			LAYER M3 ;
			RECT 80.295 254.700 80.475 254.850 ;
			LAYER M1 ;
			RECT 80.295 254.700 80.475 254.850 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[101]

	PIN QA[102]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 257.020 80.475 257.170 ;
			LAYER M2 ;
			RECT 80.295 257.020 80.475 257.170 ;
			LAYER M1 ;
			RECT 80.295 257.020 80.475 257.170 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[102]

	PIN QA[103]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 259.340 80.475 259.490 ;
			LAYER M2 ;
			RECT 80.295 259.340 80.475 259.490 ;
			LAYER M3 ;
			RECT 80.295 259.340 80.475 259.490 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[103]

	PIN QA[104]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 261.660 80.475 261.810 ;
			LAYER M2 ;
			RECT 80.295 261.660 80.475 261.810 ;
			LAYER M3 ;
			RECT 80.295 261.660 80.475 261.810 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[104]

	PIN QA[105]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 263.980 80.475 264.130 ;
			LAYER M3 ;
			RECT 80.295 263.980 80.475 264.130 ;
			LAYER M1 ;
			RECT 80.295 263.980 80.475 264.130 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[105]

	PIN QA[106]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 266.300 80.475 266.450 ;
			LAYER M1 ;
			RECT 80.295 266.300 80.475 266.450 ;
			LAYER M3 ;
			RECT 80.295 266.300 80.475 266.450 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[106]

	PIN QA[107]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 268.620 80.475 268.770 ;
			LAYER M3 ;
			RECT 80.295 268.620 80.475 268.770 ;
			LAYER M1 ;
			RECT 80.295 268.620 80.475 268.770 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[107]

	PIN QA[108]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 270.940 80.475 271.090 ;
			LAYER M1 ;
			RECT 80.295 270.940 80.475 271.090 ;
			LAYER M3 ;
			RECT 80.295 270.940 80.475 271.090 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[108]

	PIN QA[109]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 273.260 80.475 273.410 ;
			LAYER M1 ;
			RECT 80.295 273.260 80.475 273.410 ;
			LAYER M3 ;
			RECT 80.295 273.260 80.475 273.410 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[109]

	PIN QA[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 25.060 80.475 25.210 ;
			LAYER M1 ;
			RECT 80.295 25.060 80.475 25.210 ;
			LAYER M2 ;
			RECT 80.295 25.060 80.475 25.210 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[10]

	PIN QA[110]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 275.580 80.475 275.730 ;
			LAYER M1 ;
			RECT 80.295 275.580 80.475 275.730 ;
			LAYER M2 ;
			RECT 80.295 275.580 80.475 275.730 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[110]

	PIN QA[111]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 277.900 80.475 278.050 ;
			LAYER M3 ;
			RECT 80.295 277.900 80.475 278.050 ;
			LAYER M1 ;
			RECT 80.295 277.900 80.475 278.050 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[111]

	PIN QA[112]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 280.220 80.475 280.370 ;
			LAYER M3 ;
			RECT 80.295 280.220 80.475 280.370 ;
			LAYER M1 ;
			RECT 80.295 280.220 80.475 280.370 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[112]

	PIN QA[113]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 282.540 80.475 282.690 ;
			LAYER M3 ;
			RECT 80.295 282.540 80.475 282.690 ;
			LAYER M1 ;
			RECT 80.295 282.540 80.475 282.690 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[113]

	PIN QA[114]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 284.860 80.475 285.010 ;
			LAYER M1 ;
			RECT 80.295 284.860 80.475 285.010 ;
			LAYER M2 ;
			RECT 80.295 284.860 80.475 285.010 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[114]

	PIN QA[115]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 287.180 80.475 287.330 ;
			LAYER M1 ;
			RECT 80.295 287.180 80.475 287.330 ;
			LAYER M3 ;
			RECT 80.295 287.180 80.475 287.330 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[115]

	PIN QA[116]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 289.500 80.475 289.650 ;
			LAYER M3 ;
			RECT 80.295 289.500 80.475 289.650 ;
			LAYER M1 ;
			RECT 80.295 289.500 80.475 289.650 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[116]

	PIN QA[117]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 291.820 80.475 291.970 ;
			LAYER M3 ;
			RECT 80.295 291.820 80.475 291.970 ;
			LAYER M1 ;
			RECT 80.295 291.820 80.475 291.970 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[117]

	PIN QA[118]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 294.140 80.475 294.290 ;
			LAYER M3 ;
			RECT 80.295 294.140 80.475 294.290 ;
			LAYER M1 ;
			RECT 80.295 294.140 80.475 294.290 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[118]

	PIN QA[119]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 296.460 80.475 296.610 ;
			LAYER M2 ;
			RECT 80.295 296.460 80.475 296.610 ;
			LAYER M1 ;
			RECT 80.295 296.460 80.475 296.610 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[119]

	PIN QA[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 27.380 80.475 27.530 ;
			LAYER M1 ;
			RECT 80.295 27.380 80.475 27.530 ;
			LAYER M2 ;
			RECT 80.295 27.380 80.475 27.530 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[11]

	PIN QA[120]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 298.780 80.475 298.930 ;
			LAYER M2 ;
			RECT 80.295 298.780 80.475 298.930 ;
			LAYER M1 ;
			RECT 80.295 298.780 80.475 298.930 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[120]

	PIN QA[121]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 301.100 80.475 301.250 ;
			LAYER M1 ;
			RECT 80.295 301.100 80.475 301.250 ;
			LAYER M2 ;
			RECT 80.295 301.100 80.475 301.250 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[121]

	PIN QA[122]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 303.420 80.475 303.570 ;
			LAYER M3 ;
			RECT 80.295 303.420 80.475 303.570 ;
			LAYER M2 ;
			RECT 80.295 303.420 80.475 303.570 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[122]

	PIN QA[123]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 305.740 80.475 305.890 ;
			LAYER M3 ;
			RECT 80.295 305.740 80.475 305.890 ;
			LAYER M1 ;
			RECT 80.295 305.740 80.475 305.890 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[123]

	PIN QA[124]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 308.060 80.475 308.210 ;
			LAYER M2 ;
			RECT 80.295 308.060 80.475 308.210 ;
			LAYER M1 ;
			RECT 80.295 308.060 80.475 308.210 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[124]

	PIN QA[125]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 310.380 80.475 310.530 ;
			LAYER M2 ;
			RECT 80.295 310.380 80.475 310.530 ;
			LAYER M3 ;
			RECT 80.295 310.380 80.475 310.530 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[125]

	PIN QA[126]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 312.700 80.475 312.850 ;
			LAYER M1 ;
			RECT 80.295 312.700 80.475 312.850 ;
			LAYER M2 ;
			RECT 80.295 312.700 80.475 312.850 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[126]

	PIN QA[127]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 315.020 80.475 315.170 ;
			LAYER M3 ;
			RECT 80.295 315.020 80.475 315.170 ;
			LAYER M1 ;
			RECT 80.295 315.020 80.475 315.170 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[127]

	PIN QA[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 29.700 80.475 29.850 ;
			LAYER M2 ;
			RECT 80.295 29.700 80.475 29.850 ;
			LAYER M3 ;
			RECT 80.295 29.700 80.475 29.850 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[12]

	PIN QA[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 32.020 80.475 32.170 ;
			LAYER M3 ;
			RECT 80.295 32.020 80.475 32.170 ;
			LAYER M1 ;
			RECT 80.295 32.020 80.475 32.170 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[13]

	PIN QA[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 34.340 80.475 34.490 ;
			LAYER M3 ;
			RECT 80.295 34.340 80.475 34.490 ;
			LAYER M1 ;
			RECT 80.295 34.340 80.475 34.490 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[14]

	PIN QA[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 36.660 80.475 36.810 ;
			LAYER M1 ;
			RECT 80.295 36.660 80.475 36.810 ;
			LAYER M2 ;
			RECT 80.295 36.660 80.475 36.810 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[15]

	PIN QA[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 38.980 80.475 39.130 ;
			LAYER M2 ;
			RECT 80.295 38.980 80.475 39.130 ;
			LAYER M1 ;
			RECT 80.295 38.980 80.475 39.130 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[16]

	PIN QA[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 41.300 80.475 41.450 ;
			LAYER M1 ;
			RECT 80.295 41.300 80.475 41.450 ;
			LAYER M3 ;
			RECT 80.295 41.300 80.475 41.450 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[17]

	PIN QA[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 43.620 80.475 43.770 ;
			LAYER M3 ;
			RECT 80.295 43.620 80.475 43.770 ;
			LAYER M2 ;
			RECT 80.295 43.620 80.475 43.770 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[18]

	PIN QA[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 45.940 80.475 46.090 ;
			LAYER M3 ;
			RECT 80.295 45.940 80.475 46.090 ;
			LAYER M1 ;
			RECT 80.295 45.940 80.475 46.090 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[19]

	PIN QA[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 4.180 80.475 4.330 ;
			LAYER M3 ;
			RECT 80.295 4.180 80.475 4.330 ;
			LAYER M1 ;
			RECT 80.295 4.180 80.475 4.330 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[1]

	PIN QA[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 48.260 80.475 48.410 ;
			LAYER M1 ;
			RECT 80.295 48.260 80.475 48.410 ;
			LAYER M2 ;
			RECT 80.295 48.260 80.475 48.410 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[20]

	PIN QA[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 50.580 80.475 50.730 ;
			LAYER M3 ;
			RECT 80.295 50.580 80.475 50.730 ;
			LAYER M1 ;
			RECT 80.295 50.580 80.475 50.730 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[21]

	PIN QA[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 52.900 80.475 53.050 ;
			LAYER M1 ;
			RECT 80.295 52.900 80.475 53.050 ;
			LAYER M2 ;
			RECT 80.295 52.900 80.475 53.050 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[22]

	PIN QA[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 55.220 80.475 55.370 ;
			LAYER M3 ;
			RECT 80.295 55.220 80.475 55.370 ;
			LAYER M2 ;
			RECT 80.295 55.220 80.475 55.370 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[23]

	PIN QA[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 57.540 80.475 57.690 ;
			LAYER M2 ;
			RECT 80.295 57.540 80.475 57.690 ;
			LAYER M1 ;
			RECT 80.295 57.540 80.475 57.690 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[24]

	PIN QA[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 59.860 80.475 60.010 ;
			LAYER M2 ;
			RECT 80.295 59.860 80.475 60.010 ;
			LAYER M1 ;
			RECT 80.295 59.860 80.475 60.010 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[25]

	PIN QA[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 62.180 80.475 62.330 ;
			LAYER M1 ;
			RECT 80.295 62.180 80.475 62.330 ;
			LAYER M3 ;
			RECT 80.295 62.180 80.475 62.330 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[26]

	PIN QA[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 64.500 80.475 64.650 ;
			LAYER M3 ;
			RECT 80.295 64.500 80.475 64.650 ;
			LAYER M2 ;
			RECT 80.295 64.500 80.475 64.650 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[27]

	PIN QA[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 66.820 80.475 66.970 ;
			LAYER M1 ;
			RECT 80.295 66.820 80.475 66.970 ;
			LAYER M2 ;
			RECT 80.295 66.820 80.475 66.970 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[28]

	PIN QA[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 69.140 80.475 69.290 ;
			LAYER M1 ;
			RECT 80.295 69.140 80.475 69.290 ;
			LAYER M2 ;
			RECT 80.295 69.140 80.475 69.290 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[29]

	PIN QA[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 6.500 80.475 6.650 ;
			LAYER M3 ;
			RECT 80.295 6.500 80.475 6.650 ;
			LAYER M1 ;
			RECT 80.295 6.500 80.475 6.650 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[2]

	PIN QA[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 71.460 80.475 71.610 ;
			LAYER M1 ;
			RECT 80.295 71.460 80.475 71.610 ;
			LAYER M2 ;
			RECT 80.295 71.460 80.475 71.610 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[30]

	PIN QA[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 73.780 80.475 73.930 ;
			LAYER M1 ;
			RECT 80.295 73.780 80.475 73.930 ;
			LAYER M2 ;
			RECT 80.295 73.780 80.475 73.930 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[31]

	PIN QA[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 76.100 80.475 76.250 ;
			LAYER M3 ;
			RECT 80.295 76.100 80.475 76.250 ;
			LAYER M1 ;
			RECT 80.295 76.100 80.475 76.250 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[32]

	PIN QA[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 78.420 80.475 78.570 ;
			LAYER M2 ;
			RECT 80.295 78.420 80.475 78.570 ;
			LAYER M1 ;
			RECT 80.295 78.420 80.475 78.570 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[33]

	PIN QA[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 80.740 80.475 80.890 ;
			LAYER M1 ;
			RECT 80.295 80.740 80.475 80.890 ;
			LAYER M3 ;
			RECT 80.295 80.740 80.475 80.890 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[34]

	PIN QA[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 83.060 80.475 83.210 ;
			LAYER M3 ;
			RECT 80.295 83.060 80.475 83.210 ;
			LAYER M2 ;
			RECT 80.295 83.060 80.475 83.210 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[35]

	PIN QA[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 85.380 80.475 85.530 ;
			LAYER M3 ;
			RECT 80.295 85.380 80.475 85.530 ;
			LAYER M2 ;
			RECT 80.295 85.380 80.475 85.530 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[36]

	PIN QA[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 87.700 80.475 87.850 ;
			LAYER M2 ;
			RECT 80.295 87.700 80.475 87.850 ;
			LAYER M1 ;
			RECT 80.295 87.700 80.475 87.850 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[37]

	PIN QA[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 90.020 80.475 90.170 ;
			LAYER M2 ;
			RECT 80.295 90.020 80.475 90.170 ;
			LAYER M1 ;
			RECT 80.295 90.020 80.475 90.170 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[38]

	PIN QA[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 92.340 80.475 92.490 ;
			LAYER M3 ;
			RECT 80.295 92.340 80.475 92.490 ;
			LAYER M1 ;
			RECT 80.295 92.340 80.475 92.490 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[39]

	PIN QA[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 8.820 80.475 8.970 ;
			LAYER M2 ;
			RECT 80.295 8.820 80.475 8.970 ;
			LAYER M3 ;
			RECT 80.295 8.820 80.475 8.970 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[3]

	PIN QA[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 94.660 80.475 94.810 ;
			LAYER M3 ;
			RECT 80.295 94.660 80.475 94.810 ;
			LAYER M1 ;
			RECT 80.295 94.660 80.475 94.810 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[40]

	PIN QA[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 96.980 80.475 97.130 ;
			LAYER M1 ;
			RECT 80.295 96.980 80.475 97.130 ;
			LAYER M3 ;
			RECT 80.295 96.980 80.475 97.130 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[41]

	PIN QA[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 99.300 80.475 99.450 ;
			LAYER M1 ;
			RECT 80.295 99.300 80.475 99.450 ;
			LAYER M2 ;
			RECT 80.295 99.300 80.475 99.450 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[42]

	PIN QA[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 101.620 80.475 101.770 ;
			LAYER M3 ;
			RECT 80.295 101.620 80.475 101.770 ;
			LAYER M2 ;
			RECT 80.295 101.620 80.475 101.770 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[43]

	PIN QA[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 103.940 80.475 104.090 ;
			LAYER M2 ;
			RECT 80.295 103.940 80.475 104.090 ;
			LAYER M1 ;
			RECT 80.295 103.940 80.475 104.090 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[44]

	PIN QA[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 106.260 80.475 106.410 ;
			LAYER M3 ;
			RECT 80.295 106.260 80.475 106.410 ;
			LAYER M2 ;
			RECT 80.295 106.260 80.475 106.410 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[45]

	PIN QA[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 108.580 80.475 108.730 ;
			LAYER M3 ;
			RECT 80.295 108.580 80.475 108.730 ;
			LAYER M1 ;
			RECT 80.295 108.580 80.475 108.730 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[46]

	PIN QA[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 110.900 80.475 111.050 ;
			LAYER M1 ;
			RECT 80.295 110.900 80.475 111.050 ;
			LAYER M3 ;
			RECT 80.295 110.900 80.475 111.050 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[47]

	PIN QA[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 113.220 80.475 113.370 ;
			LAYER M1 ;
			RECT 80.295 113.220 80.475 113.370 ;
			LAYER M2 ;
			RECT 80.295 113.220 80.475 113.370 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[48]

	PIN QA[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 115.540 80.475 115.690 ;
			LAYER M2 ;
			RECT 80.295 115.540 80.475 115.690 ;
			LAYER M3 ;
			RECT 80.295 115.540 80.475 115.690 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[49]

	PIN QA[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 11.140 80.475 11.290 ;
			LAYER M2 ;
			RECT 80.295 11.140 80.475 11.290 ;
			LAYER M1 ;
			RECT 80.295 11.140 80.475 11.290 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[4]

	PIN QA[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 117.860 80.475 118.010 ;
			LAYER M3 ;
			RECT 80.295 117.860 80.475 118.010 ;
			LAYER M1 ;
			RECT 80.295 117.860 80.475 118.010 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[50]

	PIN QA[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 120.180 80.475 120.330 ;
			LAYER M2 ;
			RECT 80.295 120.180 80.475 120.330 ;
			LAYER M3 ;
			RECT 80.295 120.180 80.475 120.330 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[51]

	PIN QA[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 122.500 80.475 122.650 ;
			LAYER M3 ;
			RECT 80.295 122.500 80.475 122.650 ;
			LAYER M1 ;
			RECT 80.295 122.500 80.475 122.650 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[52]

	PIN QA[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 124.820 80.475 124.970 ;
			LAYER M1 ;
			RECT 80.295 124.820 80.475 124.970 ;
			LAYER M3 ;
			RECT 80.295 124.820 80.475 124.970 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[53]

	PIN QA[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 127.140 80.475 127.290 ;
			LAYER M1 ;
			RECT 80.295 127.140 80.475 127.290 ;
			LAYER M3 ;
			RECT 80.295 127.140 80.475 127.290 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[54]

	PIN QA[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 129.460 80.475 129.610 ;
			LAYER M2 ;
			RECT 80.295 129.460 80.475 129.610 ;
			LAYER M3 ;
			RECT 80.295 129.460 80.475 129.610 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[55]

	PIN QA[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 131.780 80.475 131.930 ;
			LAYER M3 ;
			RECT 80.295 131.780 80.475 131.930 ;
			LAYER M1 ;
			RECT 80.295 131.780 80.475 131.930 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[56]

	PIN QA[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 134.100 80.475 134.250 ;
			LAYER M1 ;
			RECT 80.295 134.100 80.475 134.250 ;
			LAYER M2 ;
			RECT 80.295 134.100 80.475 134.250 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[57]

	PIN QA[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 136.420 80.475 136.570 ;
			LAYER M2 ;
			RECT 80.295 136.420 80.475 136.570 ;
			LAYER M3 ;
			RECT 80.295 136.420 80.475 136.570 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[58]

	PIN QA[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 138.735 80.475 138.885 ;
			LAYER M1 ;
			RECT 80.295 138.735 80.475 138.885 ;
			LAYER M2 ;
			RECT 80.295 138.735 80.475 138.885 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[59]

	PIN QA[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 13.460 80.475 13.610 ;
			LAYER M1 ;
			RECT 80.295 13.460 80.475 13.610 ;
			LAYER M3 ;
			RECT 80.295 13.460 80.475 13.610 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[5]

	PIN QA[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 141.045 80.475 141.195 ;
			LAYER M3 ;
			RECT 80.295 141.045 80.475 141.195 ;
			LAYER M1 ;
			RECT 80.295 141.045 80.475 141.195 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[60]

	PIN QA[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 143.025 80.475 143.175 ;
			LAYER M3 ;
			RECT 80.295 143.025 80.475 143.175 ;
			LAYER M2 ;
			RECT 80.295 143.025 80.475 143.175 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[61]

	PIN QA[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 145.920 80.475 146.070 ;
			LAYER M2 ;
			RECT 80.295 145.920 80.475 146.070 ;
			LAYER M1 ;
			RECT 80.295 145.920 80.475 146.070 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[62]

	PIN QA[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 147.920 80.475 148.070 ;
			LAYER M1 ;
			RECT 80.295 147.920 80.475 148.070 ;
			LAYER M2 ;
			RECT 80.295 147.920 80.475 148.070 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[63]

	PIN QA[64]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 168.270 80.475 168.420 ;
			LAYER M3 ;
			RECT 80.295 168.270 80.475 168.420 ;
			LAYER M1 ;
			RECT 80.295 168.270 80.475 168.420 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[64]

	PIN QA[65]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 170.880 80.475 171.030 ;
			LAYER M1 ;
			RECT 80.295 170.880 80.475 171.030 ;
			LAYER M2 ;
			RECT 80.295 170.880 80.475 171.030 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[65]

	PIN QA[66]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 173.190 80.475 173.340 ;
			LAYER M1 ;
			RECT 80.295 173.190 80.475 173.340 ;
			LAYER M2 ;
			RECT 80.295 173.190 80.475 173.340 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[66]

	PIN QA[67]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 176.160 80.475 176.310 ;
			LAYER M1 ;
			RECT 80.295 176.160 80.475 176.310 ;
			LAYER M3 ;
			RECT 80.295 176.160 80.475 176.310 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[67]

	PIN QA[68]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 178.470 80.475 178.620 ;
			LAYER M3 ;
			RECT 80.295 178.470 80.475 178.620 ;
			LAYER M2 ;
			RECT 80.295 178.470 80.475 178.620 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[68]

	PIN QA[69]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 180.460 80.475 180.610 ;
			LAYER M1 ;
			RECT 80.295 180.460 80.475 180.610 ;
			LAYER M2 ;
			RECT 80.295 180.460 80.475 180.610 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[69]

	PIN QA[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 15.780 80.475 15.930 ;
			LAYER M2 ;
			RECT 80.295 15.780 80.475 15.930 ;
			LAYER M3 ;
			RECT 80.295 15.780 80.475 15.930 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[6]

	PIN QA[70]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 182.780 80.475 182.930 ;
			LAYER M1 ;
			RECT 80.295 182.780 80.475 182.930 ;
			LAYER M3 ;
			RECT 80.295 182.780 80.475 182.930 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[70]

	PIN QA[71]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 185.100 80.475 185.250 ;
			LAYER M2 ;
			RECT 80.295 185.100 80.475 185.250 ;
			LAYER M3 ;
			RECT 80.295 185.100 80.475 185.250 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[71]

	PIN QA[72]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 187.420 80.475 187.570 ;
			LAYER M2 ;
			RECT 80.295 187.420 80.475 187.570 ;
			LAYER M3 ;
			RECT 80.295 187.420 80.475 187.570 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[72]

	PIN QA[73]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 189.740 80.475 189.890 ;
			LAYER M2 ;
			RECT 80.295 189.740 80.475 189.890 ;
			LAYER M3 ;
			RECT 80.295 189.740 80.475 189.890 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[73]

	PIN QA[74]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 192.060 80.475 192.210 ;
			LAYER M1 ;
			RECT 80.295 192.060 80.475 192.210 ;
			LAYER M3 ;
			RECT 80.295 192.060 80.475 192.210 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[74]

	PIN QA[75]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 194.380 80.475 194.530 ;
			LAYER M2 ;
			RECT 80.295 194.380 80.475 194.530 ;
			LAYER M1 ;
			RECT 80.295 194.380 80.475 194.530 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[75]

	PIN QA[76]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 196.700 80.475 196.850 ;
			LAYER M2 ;
			RECT 80.295 196.700 80.475 196.850 ;
			LAYER M3 ;
			RECT 80.295 196.700 80.475 196.850 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[76]

	PIN QA[77]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 199.020 80.475 199.170 ;
			LAYER M2 ;
			RECT 80.295 199.020 80.475 199.170 ;
			LAYER M3 ;
			RECT 80.295 199.020 80.475 199.170 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[77]

	PIN QA[78]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 201.340 80.475 201.490 ;
			LAYER M1 ;
			RECT 80.295 201.340 80.475 201.490 ;
			LAYER M2 ;
			RECT 80.295 201.340 80.475 201.490 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[78]

	PIN QA[79]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 203.660 80.475 203.810 ;
			LAYER M2 ;
			RECT 80.295 203.660 80.475 203.810 ;
			LAYER M3 ;
			RECT 80.295 203.660 80.475 203.810 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[79]

	PIN QA[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 18.100 80.475 18.250 ;
			LAYER M2 ;
			RECT 80.295 18.100 80.475 18.250 ;
			LAYER M3 ;
			RECT 80.295 18.100 80.475 18.250 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[7]

	PIN QA[80]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 205.980 80.475 206.130 ;
			LAYER M3 ;
			RECT 80.295 205.980 80.475 206.130 ;
			LAYER M2 ;
			RECT 80.295 205.980 80.475 206.130 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[80]

	PIN QA[81]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 208.300 80.475 208.450 ;
			LAYER M2 ;
			RECT 80.295 208.300 80.475 208.450 ;
			LAYER M1 ;
			RECT 80.295 208.300 80.475 208.450 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[81]

	PIN QA[82]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 210.620 80.475 210.770 ;
			LAYER M3 ;
			RECT 80.295 210.620 80.475 210.770 ;
			LAYER M2 ;
			RECT 80.295 210.620 80.475 210.770 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[82]

	PIN QA[83]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 212.940 80.475 213.090 ;
			LAYER M3 ;
			RECT 80.295 212.940 80.475 213.090 ;
			LAYER M2 ;
			RECT 80.295 212.940 80.475 213.090 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[83]

	PIN QA[84]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 215.260 80.475 215.410 ;
			LAYER M1 ;
			RECT 80.295 215.260 80.475 215.410 ;
			LAYER M2 ;
			RECT 80.295 215.260 80.475 215.410 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[84]

	PIN QA[85]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 217.580 80.475 217.730 ;
			LAYER M3 ;
			RECT 80.295 217.580 80.475 217.730 ;
			LAYER M2 ;
			RECT 80.295 217.580 80.475 217.730 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[85]

	PIN QA[86]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 219.900 80.475 220.050 ;
			LAYER M3 ;
			RECT 80.295 219.900 80.475 220.050 ;
			LAYER M1 ;
			RECT 80.295 219.900 80.475 220.050 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[86]

	PIN QA[87]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 222.220 80.475 222.370 ;
			LAYER M1 ;
			RECT 80.295 222.220 80.475 222.370 ;
			LAYER M2 ;
			RECT 80.295 222.220 80.475 222.370 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[87]

	PIN QA[88]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 224.540 80.475 224.690 ;
			LAYER M1 ;
			RECT 80.295 224.540 80.475 224.690 ;
			LAYER M3 ;
			RECT 80.295 224.540 80.475 224.690 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[88]

	PIN QA[89]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 226.860 80.475 227.010 ;
			LAYER M3 ;
			RECT 80.295 226.860 80.475 227.010 ;
			LAYER M1 ;
			RECT 80.295 226.860 80.475 227.010 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[89]

	PIN QA[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 20.420 80.475 20.570 ;
			LAYER M1 ;
			RECT 80.295 20.420 80.475 20.570 ;
			LAYER M3 ;
			RECT 80.295 20.420 80.475 20.570 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[8]

	PIN QA[90]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 229.180 80.475 229.330 ;
			LAYER M3 ;
			RECT 80.295 229.180 80.475 229.330 ;
			LAYER M1 ;
			RECT 80.295 229.180 80.475 229.330 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[90]

	PIN QA[91]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 231.500 80.475 231.650 ;
			LAYER M1 ;
			RECT 80.295 231.500 80.475 231.650 ;
			LAYER M2 ;
			RECT 80.295 231.500 80.475 231.650 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[91]

	PIN QA[92]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 233.820 80.475 233.970 ;
			LAYER M3 ;
			RECT 80.295 233.820 80.475 233.970 ;
			LAYER M1 ;
			RECT 80.295 233.820 80.475 233.970 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[92]

	PIN QA[93]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 236.140 80.475 236.290 ;
			LAYER M3 ;
			RECT 80.295 236.140 80.475 236.290 ;
			LAYER M1 ;
			RECT 80.295 236.140 80.475 236.290 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[93]

	PIN QA[94]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 238.460 80.475 238.610 ;
			LAYER M3 ;
			RECT 80.295 238.460 80.475 238.610 ;
			LAYER M2 ;
			RECT 80.295 238.460 80.475 238.610 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[94]

	PIN QA[95]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 240.780 80.475 240.930 ;
			LAYER M3 ;
			RECT 80.295 240.780 80.475 240.930 ;
			LAYER M1 ;
			RECT 80.295 240.780 80.475 240.930 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[95]

	PIN QA[96]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 243.100 80.475 243.250 ;
			LAYER M1 ;
			RECT 80.295 243.100 80.475 243.250 ;
			LAYER M2 ;
			RECT 80.295 243.100 80.475 243.250 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[96]

	PIN QA[97]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 245.420 80.475 245.570 ;
			LAYER M2 ;
			RECT 80.295 245.420 80.475 245.570 ;
			LAYER M1 ;
			RECT 80.295 245.420 80.475 245.570 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[97]

	PIN QA[98]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 247.740 80.475 247.890 ;
			LAYER M3 ;
			RECT 80.295 247.740 80.475 247.890 ;
			LAYER M1 ;
			RECT 80.295 247.740 80.475 247.890 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[98]

	PIN QA[99]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 250.060 80.475 250.210 ;
			LAYER M1 ;
			RECT 80.295 250.060 80.475 250.210 ;
			LAYER M2 ;
			RECT 80.295 250.060 80.475 250.210 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[99]

	PIN QA[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 22.740 80.475 22.890 ;
			LAYER M3 ;
			RECT 80.295 22.740 80.475 22.890 ;
			LAYER M2 ;
			RECT 80.295 22.740 80.475 22.890 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[9]

	PIN QB[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 2.525 80.475 2.675 ;
			LAYER M1 ;
			RECT 80.295 2.525 80.475 2.675 ;
			LAYER M2 ;
			RECT 80.295 2.525 80.475 2.675 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[0]

	PIN QB[100]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 253.045 80.475 253.195 ;
			LAYER M2 ;
			RECT 80.295 253.045 80.475 253.195 ;
			LAYER M1 ;
			RECT 80.295 253.045 80.475 253.195 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[100]

	PIN QB[101]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 255.365 80.475 255.515 ;
			LAYER M2 ;
			RECT 80.295 255.365 80.475 255.515 ;
			LAYER M1 ;
			RECT 80.295 255.365 80.475 255.515 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[101]

	PIN QB[102]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 257.685 80.475 257.835 ;
			LAYER M1 ;
			RECT 80.295 257.685 80.475 257.835 ;
			LAYER M2 ;
			RECT 80.295 257.685 80.475 257.835 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[102]

	PIN QB[103]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 260.005 80.475 260.155 ;
			LAYER M1 ;
			RECT 80.295 260.005 80.475 260.155 ;
			LAYER M2 ;
			RECT 80.295 260.005 80.475 260.155 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[103]

	PIN QB[104]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 262.325 80.475 262.475 ;
			LAYER M1 ;
			RECT 80.295 262.325 80.475 262.475 ;
			LAYER M3 ;
			RECT 80.295 262.325 80.475 262.475 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[104]

	PIN QB[105]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 264.645 80.475 264.795 ;
			LAYER M1 ;
			RECT 80.295 264.645 80.475 264.795 ;
			LAYER M2 ;
			RECT 80.295 264.645 80.475 264.795 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[105]

	PIN QB[106]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 266.965 80.475 267.115 ;
			LAYER M3 ;
			RECT 80.295 266.965 80.475 267.115 ;
			LAYER M2 ;
			RECT 80.295 266.965 80.475 267.115 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[106]

	PIN QB[107]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 269.285 80.475 269.435 ;
			LAYER M1 ;
			RECT 80.295 269.285 80.475 269.435 ;
			LAYER M3 ;
			RECT 80.295 269.285 80.475 269.435 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[107]

	PIN QB[108]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 271.605 80.475 271.755 ;
			LAYER M2 ;
			RECT 80.295 271.605 80.475 271.755 ;
			LAYER M1 ;
			RECT 80.295 271.605 80.475 271.755 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[108]

	PIN QB[109]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 273.925 80.475 274.075 ;
			LAYER M1 ;
			RECT 80.295 273.925 80.475 274.075 ;
			LAYER M2 ;
			RECT 80.295 273.925 80.475 274.075 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[109]

	PIN QB[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 25.725 80.475 25.875 ;
			LAYER M1 ;
			RECT 80.295 25.725 80.475 25.875 ;
			LAYER M2 ;
			RECT 80.295 25.725 80.475 25.875 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[10]

	PIN QB[110]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 276.245 80.475 276.395 ;
			LAYER M3 ;
			RECT 80.295 276.245 80.475 276.395 ;
			LAYER M1 ;
			RECT 80.295 276.245 80.475 276.395 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[110]

	PIN QB[111]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 278.565 80.475 278.715 ;
			LAYER M1 ;
			RECT 80.295 278.565 80.475 278.715 ;
			LAYER M2 ;
			RECT 80.295 278.565 80.475 278.715 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[111]

	PIN QB[112]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 280.885 80.475 281.035 ;
			LAYER M3 ;
			RECT 80.295 280.885 80.475 281.035 ;
			LAYER M1 ;
			RECT 80.295 280.885 80.475 281.035 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[112]

	PIN QB[113]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 283.205 80.475 283.355 ;
			LAYER M1 ;
			RECT 80.295 283.205 80.475 283.355 ;
			LAYER M2 ;
			RECT 80.295 283.205 80.475 283.355 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[113]

	PIN QB[114]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 285.525 80.475 285.675 ;
			LAYER M2 ;
			RECT 80.295 285.525 80.475 285.675 ;
			LAYER M1 ;
			RECT 80.295 285.525 80.475 285.675 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[114]

	PIN QB[115]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 287.845 80.475 287.995 ;
			LAYER M1 ;
			RECT 80.295 287.845 80.475 287.995 ;
			LAYER M2 ;
			RECT 80.295 287.845 80.475 287.995 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[115]

	PIN QB[116]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 290.165 80.475 290.315 ;
			LAYER M2 ;
			RECT 80.295 290.165 80.475 290.315 ;
			LAYER M1 ;
			RECT 80.295 290.165 80.475 290.315 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[116]

	PIN QB[117]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 292.485 80.475 292.635 ;
			LAYER M2 ;
			RECT 80.295 292.485 80.475 292.635 ;
			LAYER M1 ;
			RECT 80.295 292.485 80.475 292.635 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[117]

	PIN QB[118]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 294.805 80.475 294.955 ;
			LAYER M2 ;
			RECT 80.295 294.805 80.475 294.955 ;
			LAYER M3 ;
			RECT 80.295 294.805 80.475 294.955 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[118]

	PIN QB[119]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 297.125 80.475 297.275 ;
			LAYER M1 ;
			RECT 80.295 297.125 80.475 297.275 ;
			LAYER M3 ;
			RECT 80.295 297.125 80.475 297.275 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[119]

	PIN QB[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 28.045 80.475 28.195 ;
			LAYER M3 ;
			RECT 80.295 28.045 80.475 28.195 ;
			LAYER M1 ;
			RECT 80.295 28.045 80.475 28.195 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[11]

	PIN QB[120]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 299.445 80.475 299.595 ;
			LAYER M1 ;
			RECT 80.295 299.445 80.475 299.595 ;
			LAYER M2 ;
			RECT 80.295 299.445 80.475 299.595 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[120]

	PIN QB[121]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 301.765 80.475 301.915 ;
			LAYER M1 ;
			RECT 80.295 301.765 80.475 301.915 ;
			LAYER M2 ;
			RECT 80.295 301.765 80.475 301.915 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[121]

	PIN QB[122]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 304.085 80.475 304.235 ;
			LAYER M3 ;
			RECT 80.295 304.085 80.475 304.235 ;
			LAYER M2 ;
			RECT 80.295 304.085 80.475 304.235 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[122]

	PIN QB[123]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 306.405 80.475 306.555 ;
			LAYER M3 ;
			RECT 80.295 306.405 80.475 306.555 ;
			LAYER M1 ;
			RECT 80.295 306.405 80.475 306.555 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[123]

	PIN QB[124]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 308.725 80.475 308.875 ;
			LAYER M2 ;
			RECT 80.295 308.725 80.475 308.875 ;
			LAYER M3 ;
			RECT 80.295 308.725 80.475 308.875 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[124]

	PIN QB[125]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 311.045 80.475 311.195 ;
			LAYER M1 ;
			RECT 80.295 311.045 80.475 311.195 ;
			LAYER M2 ;
			RECT 80.295 311.045 80.475 311.195 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[125]

	PIN QB[126]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 313.365 80.475 313.515 ;
			LAYER M1 ;
			RECT 80.295 313.365 80.475 313.515 ;
			LAYER M2 ;
			RECT 80.295 313.365 80.475 313.515 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[126]

	PIN QB[127]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 315.685 80.475 315.835 ;
			LAYER M1 ;
			RECT 80.295 315.685 80.475 315.835 ;
			LAYER M2 ;
			RECT 80.295 315.685 80.475 315.835 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[127]

	PIN QB[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 30.365 80.475 30.515 ;
			LAYER M2 ;
			RECT 80.295 30.365 80.475 30.515 ;
			LAYER M1 ;
			RECT 80.295 30.365 80.475 30.515 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[12]

	PIN QB[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 32.685 80.475 32.835 ;
			LAYER M3 ;
			RECT 80.295 32.685 80.475 32.835 ;
			LAYER M2 ;
			RECT 80.295 32.685 80.475 32.835 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[13]

	PIN QB[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 35.005 80.475 35.155 ;
			LAYER M3 ;
			RECT 80.295 35.005 80.475 35.155 ;
			LAYER M2 ;
			RECT 80.295 35.005 80.475 35.155 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[14]

	PIN QB[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 37.325 80.475 37.475 ;
			LAYER M2 ;
			RECT 80.295 37.325 80.475 37.475 ;
			LAYER M1 ;
			RECT 80.295 37.325 80.475 37.475 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[15]

	PIN QB[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 39.645 80.475 39.795 ;
			LAYER M2 ;
			RECT 80.295 39.645 80.475 39.795 ;
			LAYER M3 ;
			RECT 80.295 39.645 80.475 39.795 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[16]

	PIN QB[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 41.965 80.475 42.115 ;
			LAYER M2 ;
			RECT 80.295 41.965 80.475 42.115 ;
			LAYER M1 ;
			RECT 80.295 41.965 80.475 42.115 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[17]

	PIN QB[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 44.285 80.475 44.435 ;
			LAYER M1 ;
			RECT 80.295 44.285 80.475 44.435 ;
			LAYER M3 ;
			RECT 80.295 44.285 80.475 44.435 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[18]

	PIN QB[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 46.605 80.475 46.755 ;
			LAYER M2 ;
			RECT 80.295 46.605 80.475 46.755 ;
			LAYER M3 ;
			RECT 80.295 46.605 80.475 46.755 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[19]

	PIN QB[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 4.845 80.475 4.995 ;
			LAYER M3 ;
			RECT 80.295 4.845 80.475 4.995 ;
			LAYER M1 ;
			RECT 80.295 4.845 80.475 4.995 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[1]

	PIN QB[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 48.925 80.475 49.075 ;
			LAYER M1 ;
			RECT 80.295 48.925 80.475 49.075 ;
			LAYER M3 ;
			RECT 80.295 48.925 80.475 49.075 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[20]

	PIN QB[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 51.245 80.475 51.395 ;
			LAYER M2 ;
			RECT 80.295 51.245 80.475 51.395 ;
			LAYER M3 ;
			RECT 80.295 51.245 80.475 51.395 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[21]

	PIN QB[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 53.565 80.475 53.715 ;
			LAYER M2 ;
			RECT 80.295 53.565 80.475 53.715 ;
			LAYER M3 ;
			RECT 80.295 53.565 80.475 53.715 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[22]

	PIN QB[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 55.885 80.475 56.035 ;
			LAYER M3 ;
			RECT 80.295 55.885 80.475 56.035 ;
			LAYER M2 ;
			RECT 80.295 55.885 80.475 56.035 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[23]

	PIN QB[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 58.205 80.475 58.355 ;
			LAYER M2 ;
			RECT 80.295 58.205 80.475 58.355 ;
			LAYER M3 ;
			RECT 80.295 58.205 80.475 58.355 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[24]

	PIN QB[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 60.525 80.475 60.675 ;
			LAYER M3 ;
			RECT 80.295 60.525 80.475 60.675 ;
			LAYER M1 ;
			RECT 80.295 60.525 80.475 60.675 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[25]

	PIN QB[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 62.845 80.475 62.995 ;
			LAYER M2 ;
			RECT 80.295 62.845 80.475 62.995 ;
			LAYER M1 ;
			RECT 80.295 62.845 80.475 62.995 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[26]

	PIN QB[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 65.165 80.475 65.315 ;
			LAYER M3 ;
			RECT 80.295 65.165 80.475 65.315 ;
			LAYER M2 ;
			RECT 80.295 65.165 80.475 65.315 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[27]

	PIN QB[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 67.485 80.475 67.635 ;
			LAYER M2 ;
			RECT 80.295 67.485 80.475 67.635 ;
			LAYER M1 ;
			RECT 80.295 67.485 80.475 67.635 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[28]

	PIN QB[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 69.805 80.475 69.955 ;
			LAYER M1 ;
			RECT 80.295 69.805 80.475 69.955 ;
			LAYER M3 ;
			RECT 80.295 69.805 80.475 69.955 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[29]

	PIN QB[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 7.165 80.475 7.315 ;
			LAYER M2 ;
			RECT 80.295 7.165 80.475 7.315 ;
			LAYER M3 ;
			RECT 80.295 7.165 80.475 7.315 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[2]

	PIN QB[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 72.125 80.475 72.275 ;
			LAYER M3 ;
			RECT 80.295 72.125 80.475 72.275 ;
			LAYER M2 ;
			RECT 80.295 72.125 80.475 72.275 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[30]

	PIN QB[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 74.445 80.475 74.595 ;
			LAYER M2 ;
			RECT 80.295 74.445 80.475 74.595 ;
			LAYER M3 ;
			RECT 80.295 74.445 80.475 74.595 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[31]

	PIN QB[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 76.765 80.475 76.915 ;
			LAYER M1 ;
			RECT 80.295 76.765 80.475 76.915 ;
			LAYER M2 ;
			RECT 80.295 76.765 80.475 76.915 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[32]

	PIN QB[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 79.085 80.475 79.235 ;
			LAYER M2 ;
			RECT 80.295 79.085 80.475 79.235 ;
			LAYER M1 ;
			RECT 80.295 79.085 80.475 79.235 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[33]

	PIN QB[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 81.405 80.475 81.555 ;
			LAYER M1 ;
			RECT 80.295 81.405 80.475 81.555 ;
			LAYER M2 ;
			RECT 80.295 81.405 80.475 81.555 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[34]

	PIN QB[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 83.725 80.475 83.875 ;
			LAYER M3 ;
			RECT 80.295 83.725 80.475 83.875 ;
			LAYER M2 ;
			RECT 80.295 83.725 80.475 83.875 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[35]

	PIN QB[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 86.045 80.475 86.195 ;
			LAYER M2 ;
			RECT 80.295 86.045 80.475 86.195 ;
			LAYER M3 ;
			RECT 80.295 86.045 80.475 86.195 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[36]

	PIN QB[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 88.365 80.475 88.515 ;
			LAYER M1 ;
			RECT 80.295 88.365 80.475 88.515 ;
			LAYER M2 ;
			RECT 80.295 88.365 80.475 88.515 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[37]

	PIN QB[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 90.685 80.475 90.835 ;
			LAYER M1 ;
			RECT 80.295 90.685 80.475 90.835 ;
			LAYER M2 ;
			RECT 80.295 90.685 80.475 90.835 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[38]

	PIN QB[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 93.005 80.475 93.155 ;
			LAYER M1 ;
			RECT 80.295 93.005 80.475 93.155 ;
			LAYER M2 ;
			RECT 80.295 93.005 80.475 93.155 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[39]

	PIN QB[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 9.485 80.475 9.635 ;
			LAYER M2 ;
			RECT 80.295 9.485 80.475 9.635 ;
			LAYER M3 ;
			RECT 80.295 9.485 80.475 9.635 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[3]

	PIN QB[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 95.325 80.475 95.475 ;
			LAYER M1 ;
			RECT 80.295 95.325 80.475 95.475 ;
			LAYER M2 ;
			RECT 80.295 95.325 80.475 95.475 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[40]

	PIN QB[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 97.645 80.475 97.795 ;
			LAYER M1 ;
			RECT 80.295 97.645 80.475 97.795 ;
			LAYER M2 ;
			RECT 80.295 97.645 80.475 97.795 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[41]

	PIN QB[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 99.965 80.475 100.115 ;
			LAYER M1 ;
			RECT 80.295 99.965 80.475 100.115 ;
			LAYER M2 ;
			RECT 80.295 99.965 80.475 100.115 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[42]

	PIN QB[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 102.285 80.475 102.435 ;
			LAYER M3 ;
			RECT 80.295 102.285 80.475 102.435 ;
			LAYER M1 ;
			RECT 80.295 102.285 80.475 102.435 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[43]

	PIN QB[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 104.605 80.475 104.755 ;
			LAYER M1 ;
			RECT 80.295 104.605 80.475 104.755 ;
			LAYER M2 ;
			RECT 80.295 104.605 80.475 104.755 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[44]

	PIN QB[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 106.925 80.475 107.075 ;
			LAYER M1 ;
			RECT 80.295 106.925 80.475 107.075 ;
			LAYER M3 ;
			RECT 80.295 106.925 80.475 107.075 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[45]

	PIN QB[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 109.245 80.475 109.395 ;
			LAYER M1 ;
			RECT 80.295 109.245 80.475 109.395 ;
			LAYER M2 ;
			RECT 80.295 109.245 80.475 109.395 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[46]

	PIN QB[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 111.565 80.475 111.715 ;
			LAYER M2 ;
			RECT 80.295 111.565 80.475 111.715 ;
			LAYER M1 ;
			RECT 80.295 111.565 80.475 111.715 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[47]

	PIN QB[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 113.885 80.475 114.035 ;
			LAYER M2 ;
			RECT 80.295 113.885 80.475 114.035 ;
			LAYER M3 ;
			RECT 80.295 113.885 80.475 114.035 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[48]

	PIN QB[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 116.205 80.475 116.355 ;
			LAYER M1 ;
			RECT 80.295 116.205 80.475 116.355 ;
			LAYER M2 ;
			RECT 80.295 116.205 80.475 116.355 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[49]

	PIN QB[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 11.805 80.475 11.955 ;
			LAYER M2 ;
			RECT 80.295 11.805 80.475 11.955 ;
			LAYER M3 ;
			RECT 80.295 11.805 80.475 11.955 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[4]

	PIN QB[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 118.525 80.475 118.675 ;
			LAYER M2 ;
			RECT 80.295 118.525 80.475 118.675 ;
			LAYER M1 ;
			RECT 80.295 118.525 80.475 118.675 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[50]

	PIN QB[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 120.845 80.475 120.995 ;
			LAYER M2 ;
			RECT 80.295 120.845 80.475 120.995 ;
			LAYER M3 ;
			RECT 80.295 120.845 80.475 120.995 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[51]

	PIN QB[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 123.165 80.475 123.315 ;
			LAYER M1 ;
			RECT 80.295 123.165 80.475 123.315 ;
			LAYER M2 ;
			RECT 80.295 123.165 80.475 123.315 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[52]

	PIN QB[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 125.485 80.475 125.635 ;
			LAYER M1 ;
			RECT 80.295 125.485 80.475 125.635 ;
			LAYER M2 ;
			RECT 80.295 125.485 80.475 125.635 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[53]

	PIN QB[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 127.805 80.475 127.955 ;
			LAYER M3 ;
			RECT 80.295 127.805 80.475 127.955 ;
			LAYER M2 ;
			RECT 80.295 127.805 80.475 127.955 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[54]

	PIN QB[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 130.125 80.475 130.275 ;
			LAYER M2 ;
			RECT 80.295 130.125 80.475 130.275 ;
			LAYER M1 ;
			RECT 80.295 130.125 80.475 130.275 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[55]

	PIN QB[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 132.445 80.475 132.595 ;
			LAYER M1 ;
			RECT 80.295 132.445 80.475 132.595 ;
			LAYER M2 ;
			RECT 80.295 132.445 80.475 132.595 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[56]

	PIN QB[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 134.765 80.475 134.915 ;
			LAYER M2 ;
			RECT 80.295 134.765 80.475 134.915 ;
			LAYER M1 ;
			RECT 80.295 134.765 80.475 134.915 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[57]

	PIN QB[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 137.085 80.475 137.235 ;
			LAYER M1 ;
			RECT 80.295 137.085 80.475 137.235 ;
			LAYER M2 ;
			RECT 80.295 137.085 80.475 137.235 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[58]

	PIN QB[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 139.065 80.475 139.215 ;
			LAYER M2 ;
			RECT 80.295 139.065 80.475 139.215 ;
			LAYER M3 ;
			RECT 80.295 139.065 80.475 139.215 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[59]

	PIN QB[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 14.125 80.475 14.275 ;
			LAYER M1 ;
			RECT 80.295 14.125 80.475 14.275 ;
			LAYER M2 ;
			RECT 80.295 14.125 80.475 14.275 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[5]

	PIN QB[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 141.375 80.475 141.525 ;
			LAYER M2 ;
			RECT 80.295 141.375 80.475 141.525 ;
			LAYER M1 ;
			RECT 80.295 141.375 80.475 141.525 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[60]

	PIN QB[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 143.355 80.475 143.505 ;
			LAYER M1 ;
			RECT 80.295 143.355 80.475 143.505 ;
			LAYER M3 ;
			RECT 80.295 143.355 80.475 143.505 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[61]

	PIN QB[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 146.250 80.475 146.400 ;
			LAYER M3 ;
			RECT 80.295 146.250 80.475 146.400 ;
			LAYER M2 ;
			RECT 80.295 146.250 80.475 146.400 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[62]

	PIN QB[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 148.295 80.475 148.445 ;
			LAYER M2 ;
			RECT 80.295 148.295 80.475 148.445 ;
			LAYER M1 ;
			RECT 80.295 148.295 80.475 148.445 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[63]

	PIN QB[64]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 168.600 80.475 168.750 ;
			LAYER M2 ;
			RECT 80.295 168.600 80.475 168.750 ;
			LAYER M1 ;
			RECT 80.295 168.600 80.475 168.750 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[64]

	PIN QB[65]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 171.210 80.475 171.360 ;
			LAYER M2 ;
			RECT 80.295 171.210 80.475 171.360 ;
			LAYER M1 ;
			RECT 80.295 171.210 80.475 171.360 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[65]

	PIN QB[66]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 174.510 80.475 174.660 ;
			LAYER M1 ;
			RECT 80.295 174.510 80.475 174.660 ;
			LAYER M2 ;
			RECT 80.295 174.510 80.475 174.660 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[66]

	PIN QB[67]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 176.490 80.475 176.640 ;
			LAYER M3 ;
			RECT 80.295 176.490 80.475 176.640 ;
			LAYER M1 ;
			RECT 80.295 176.490 80.475 176.640 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[67]

	PIN QB[68]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 178.805 80.475 178.955 ;
			LAYER M1 ;
			RECT 80.295 178.805 80.475 178.955 ;
			LAYER M2 ;
			RECT 80.295 178.805 80.475 178.955 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[68]

	PIN QB[69]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 181.125 80.475 181.275 ;
			LAYER M2 ;
			RECT 80.295 181.125 80.475 181.275 ;
			LAYER M1 ;
			RECT 80.295 181.125 80.475 181.275 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[69]

	PIN QB[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 16.445 80.475 16.595 ;
			LAYER M1 ;
			RECT 80.295 16.445 80.475 16.595 ;
			LAYER M2 ;
			RECT 80.295 16.445 80.475 16.595 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[6]

	PIN QB[70]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 183.445 80.475 183.595 ;
			LAYER M1 ;
			RECT 80.295 183.445 80.475 183.595 ;
			LAYER M3 ;
			RECT 80.295 183.445 80.475 183.595 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[70]

	PIN QB[71]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 185.765 80.475 185.915 ;
			LAYER M3 ;
			RECT 80.295 185.765 80.475 185.915 ;
			LAYER M1 ;
			RECT 80.295 185.765 80.475 185.915 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[71]

	PIN QB[72]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 188.085 80.475 188.235 ;
			LAYER M1 ;
			RECT 80.295 188.085 80.475 188.235 ;
			LAYER M3 ;
			RECT 80.295 188.085 80.475 188.235 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[72]

	PIN QB[73]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 190.405 80.475 190.555 ;
			LAYER M2 ;
			RECT 80.295 190.405 80.475 190.555 ;
			LAYER M3 ;
			RECT 80.295 190.405 80.475 190.555 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[73]

	PIN QB[74]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 192.725 80.475 192.875 ;
			LAYER M1 ;
			RECT 80.295 192.725 80.475 192.875 ;
			LAYER M2 ;
			RECT 80.295 192.725 80.475 192.875 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[74]

	PIN QB[75]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 195.045 80.475 195.195 ;
			LAYER M1 ;
			RECT 80.295 195.045 80.475 195.195 ;
			LAYER M2 ;
			RECT 80.295 195.045 80.475 195.195 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[75]

	PIN QB[76]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 197.365 80.475 197.515 ;
			LAYER M1 ;
			RECT 80.295 197.365 80.475 197.515 ;
			LAYER M2 ;
			RECT 80.295 197.365 80.475 197.515 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[76]

	PIN QB[77]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 199.685 80.475 199.835 ;
			LAYER M3 ;
			RECT 80.295 199.685 80.475 199.835 ;
			LAYER M2 ;
			RECT 80.295 199.685 80.475 199.835 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[77]

	PIN QB[78]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 202.005 80.475 202.155 ;
			LAYER M1 ;
			RECT 80.295 202.005 80.475 202.155 ;
			LAYER M2 ;
			RECT 80.295 202.005 80.475 202.155 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[78]

	PIN QB[79]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 204.325 80.475 204.475 ;
			LAYER M2 ;
			RECT 80.295 204.325 80.475 204.475 ;
			LAYER M1 ;
			RECT 80.295 204.325 80.475 204.475 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[79]

	PIN QB[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 18.765 80.475 18.915 ;
			LAYER M1 ;
			RECT 80.295 18.765 80.475 18.915 ;
			LAYER M2 ;
			RECT 80.295 18.765 80.475 18.915 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[7]

	PIN QB[80]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 206.645 80.475 206.795 ;
			LAYER M1 ;
			RECT 80.295 206.645 80.475 206.795 ;
			LAYER M2 ;
			RECT 80.295 206.645 80.475 206.795 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[80]

	PIN QB[81]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 208.965 80.475 209.115 ;
			LAYER M1 ;
			RECT 80.295 208.965 80.475 209.115 ;
			LAYER M2 ;
			RECT 80.295 208.965 80.475 209.115 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[81]

	PIN QB[82]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 211.285 80.475 211.435 ;
			LAYER M2 ;
			RECT 80.295 211.285 80.475 211.435 ;
			LAYER M3 ;
			RECT 80.295 211.285 80.475 211.435 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[82]

	PIN QB[83]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 213.605 80.475 213.755 ;
			LAYER M3 ;
			RECT 80.295 213.605 80.475 213.755 ;
			LAYER M1 ;
			RECT 80.295 213.605 80.475 213.755 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[83]

	PIN QB[84]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 215.925 80.475 216.075 ;
			LAYER M1 ;
			RECT 80.295 215.925 80.475 216.075 ;
			LAYER M2 ;
			RECT 80.295 215.925 80.475 216.075 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[84]

	PIN QB[85]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 218.245 80.475 218.395 ;
			LAYER M3 ;
			RECT 80.295 218.245 80.475 218.395 ;
			LAYER M2 ;
			RECT 80.295 218.245 80.475 218.395 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[85]

	PIN QB[86]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 220.565 80.475 220.715 ;
			LAYER M1 ;
			RECT 80.295 220.565 80.475 220.715 ;
			LAYER M2 ;
			RECT 80.295 220.565 80.475 220.715 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[86]

	PIN QB[87]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 222.885 80.475 223.035 ;
			LAYER M1 ;
			RECT 80.295 222.885 80.475 223.035 ;
			LAYER M2 ;
			RECT 80.295 222.885 80.475 223.035 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[87]

	PIN QB[88]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 225.205 80.475 225.355 ;
			LAYER M2 ;
			RECT 80.295 225.205 80.475 225.355 ;
			LAYER M3 ;
			RECT 80.295 225.205 80.475 225.355 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[88]

	PIN QB[89]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 227.525 80.475 227.675 ;
			LAYER M3 ;
			RECT 80.295 227.525 80.475 227.675 ;
			LAYER M2 ;
			RECT 80.295 227.525 80.475 227.675 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[89]

	PIN QB[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 21.085 80.475 21.235 ;
			LAYER M2 ;
			RECT 80.295 21.085 80.475 21.235 ;
			LAYER M3 ;
			RECT 80.295 21.085 80.475 21.235 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[8]

	PIN QB[90]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 229.845 80.475 229.995 ;
			LAYER M3 ;
			RECT 80.295 229.845 80.475 229.995 ;
			LAYER M2 ;
			RECT 80.295 229.845 80.475 229.995 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[90]

	PIN QB[91]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 232.165 80.475 232.315 ;
			LAYER M2 ;
			RECT 80.295 232.165 80.475 232.315 ;
			LAYER M1 ;
			RECT 80.295 232.165 80.475 232.315 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[91]

	PIN QB[92]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 234.485 80.475 234.635 ;
			LAYER M1 ;
			RECT 80.295 234.485 80.475 234.635 ;
			LAYER M2 ;
			RECT 80.295 234.485 80.475 234.635 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[92]

	PIN QB[93]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 236.805 80.475 236.955 ;
			LAYER M1 ;
			RECT 80.295 236.805 80.475 236.955 ;
			LAYER M2 ;
			RECT 80.295 236.805 80.475 236.955 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[93]

	PIN QB[94]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 239.125 80.475 239.275 ;
			LAYER M3 ;
			RECT 80.295 239.125 80.475 239.275 ;
			LAYER M2 ;
			RECT 80.295 239.125 80.475 239.275 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[94]

	PIN QB[95]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 241.445 80.475 241.595 ;
			LAYER M3 ;
			RECT 80.295 241.445 80.475 241.595 ;
			LAYER M1 ;
			RECT 80.295 241.445 80.475 241.595 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[95]

	PIN QB[96]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 243.765 80.475 243.915 ;
			LAYER M1 ;
			RECT 80.295 243.765 80.475 243.915 ;
			LAYER M2 ;
			RECT 80.295 243.765 80.475 243.915 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[96]

	PIN QB[97]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 246.085 80.475 246.235 ;
			LAYER M1 ;
			RECT 80.295 246.085 80.475 246.235 ;
			LAYER M2 ;
			RECT 80.295 246.085 80.475 246.235 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[97]

	PIN QB[98]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 248.405 80.475 248.555 ;
			LAYER M2 ;
			RECT 80.295 248.405 80.475 248.555 ;
			LAYER M1 ;
			RECT 80.295 248.405 80.475 248.555 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[98]

	PIN QB[99]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 250.725 80.475 250.875 ;
			LAYER M2 ;
			RECT 80.295 250.725 80.475 250.875 ;
			LAYER M1 ;
			RECT 80.295 250.725 80.475 250.875 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[99]

	PIN QB[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 23.405 80.475 23.555 ;
			LAYER M1 ;
			RECT 80.295 23.405 80.475 23.555 ;
			LAYER M2 ;
			RECT 80.295 23.405 80.475 23.555 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[9]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.295 173.850 80.475 174.000 ;
			LAYER M2 ;
			RECT 80.295 173.850 80.475 174.000 ;
			LAYER M3 ;
			RECT 80.295 173.850 80.475 174.000 ;
		END
		ANTENNAGATEAREA 0.045600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.275900 LAYER M1 ;
		ANTENNAMAXAREACAR 7.227300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.393900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.045600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.199800 LAYER M2 ;
		ANTENNAMAXAREACAR 11.181800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.787900 LAYER VIA2 ;
		ANTENNAGATEAREA 0.045600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.090400 LAYER M3 ;
		ANTENNAMAXAREACAR 12.818200 LAYER M3 ;
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 174.180 80.475 174.330 ;
			LAYER M1 ;
			RECT 80.295 174.180 80.475 174.330 ;
			LAYER M2 ;
			RECT 80.295 174.180 80.475 174.330 ;
		END
		ANTENNAGATEAREA 0.045600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.275900 LAYER M1 ;
		ANTENNAMAXAREACAR 7.227300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.393900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.045600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.199800 LAYER M2 ;
		ANTENNAMAXAREACAR 11.181800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.787900 LAYER VIA2 ;
		ANTENNAGATEAREA 0.045600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.090400 LAYER M3 ;
		ANTENNAMAXAREACAR 12.818200 LAYER M3 ;
	END RTSEL[1]

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.000 1.395 80.085 1.725 ;
			LAYER M4 ;
			RECT 0.000 3.715 80.085 4.045 ;
			LAYER M4 ;
			RECT 0.000 6.035 80.085 6.365 ;
			LAYER M4 ;
			RECT 0.000 8.355 80.085 8.685 ;
			LAYER M4 ;
			RECT 0.000 10.675 80.085 11.005 ;
			LAYER M4 ;
			RECT 0.000 12.995 80.085 13.325 ;
			LAYER M4 ;
			RECT 0.000 15.315 80.085 15.645 ;
			LAYER M4 ;
			RECT 0.000 17.635 80.085 17.965 ;
			LAYER M4 ;
			RECT 0.000 19.955 80.085 20.285 ;
			LAYER M4 ;
			RECT 0.000 22.275 80.085 22.605 ;
			LAYER M4 ;
			RECT 0.000 24.595 80.085 24.925 ;
			LAYER M4 ;
			RECT 0.000 26.915 80.085 27.245 ;
			LAYER M4 ;
			RECT 0.000 29.235 80.085 29.565 ;
			LAYER M4 ;
			RECT 0.000 31.555 80.085 31.885 ;
			LAYER M4 ;
			RECT 0.000 33.875 80.085 34.205 ;
			LAYER M4 ;
			RECT 0.000 36.195 80.085 36.525 ;
			LAYER M4 ;
			RECT 0.000 38.515 80.085 38.845 ;
			LAYER M4 ;
			RECT 0.000 40.835 80.085 41.165 ;
			LAYER M4 ;
			RECT 0.000 43.155 80.085 43.485 ;
			LAYER M4 ;
			RECT 0.000 45.475 80.085 45.805 ;
			LAYER M4 ;
			RECT 0.000 47.795 80.085 48.125 ;
			LAYER M4 ;
			RECT 0.000 50.115 80.085 50.445 ;
			LAYER M4 ;
			RECT 0.000 52.435 80.085 52.765 ;
			LAYER M4 ;
			RECT 0.000 54.755 80.085 55.085 ;
			LAYER M4 ;
			RECT 0.000 57.075 80.085 57.405 ;
			LAYER M4 ;
			RECT 0.000 59.395 80.085 59.725 ;
			LAYER M4 ;
			RECT 0.000 61.715 80.085 62.045 ;
			LAYER M4 ;
			RECT 0.000 64.035 80.085 64.365 ;
			LAYER M4 ;
			RECT 0.000 66.355 80.085 66.685 ;
			LAYER M4 ;
			RECT 0.000 68.675 80.085 69.005 ;
			LAYER M4 ;
			RECT 0.000 70.995 80.085 71.325 ;
			LAYER M4 ;
			RECT 0.000 73.315 80.085 73.645 ;
			LAYER M4 ;
			RECT 0.000 75.635 80.085 75.965 ;
			LAYER M4 ;
			RECT 0.000 77.955 80.085 78.285 ;
			LAYER M4 ;
			RECT 0.000 80.275 80.085 80.605 ;
			LAYER M4 ;
			RECT 0.000 82.595 80.085 82.925 ;
			LAYER M4 ;
			RECT 0.000 84.915 80.085 85.245 ;
			LAYER M4 ;
			RECT 0.000 87.235 80.085 87.565 ;
			LAYER M4 ;
			RECT 0.000 89.555 80.085 89.885 ;
			LAYER M4 ;
			RECT 0.000 91.875 80.085 92.205 ;
			LAYER M4 ;
			RECT 0.000 94.195 80.085 94.525 ;
			LAYER M4 ;
			RECT 0.000 96.515 80.085 96.845 ;
			LAYER M4 ;
			RECT 0.000 98.835 80.085 99.165 ;
			LAYER M4 ;
			RECT 0.000 101.155 80.085 101.485 ;
			LAYER M4 ;
			RECT 0.000 103.475 80.085 103.805 ;
			LAYER M4 ;
			RECT 0.000 105.795 80.085 106.125 ;
			LAYER M4 ;
			RECT 0.000 108.115 80.085 108.445 ;
			LAYER M4 ;
			RECT 0.000 110.435 80.085 110.765 ;
			LAYER M4 ;
			RECT 0.000 112.755 80.085 113.085 ;
			LAYER M4 ;
			RECT 0.000 115.075 80.085 115.405 ;
			LAYER M4 ;
			RECT 0.000 117.395 80.085 117.725 ;
			LAYER M4 ;
			RECT 0.000 119.715 80.085 120.045 ;
			LAYER M4 ;
			RECT 0.000 122.035 80.085 122.365 ;
			LAYER M4 ;
			RECT 0.000 124.355 80.085 124.685 ;
			LAYER M4 ;
			RECT 0.000 126.675 80.085 127.005 ;
			LAYER M4 ;
			RECT 0.000 128.995 80.085 129.325 ;
			LAYER M4 ;
			RECT 0.000 131.315 80.085 131.645 ;
			LAYER M4 ;
			RECT 0.000 133.635 80.085 133.965 ;
			LAYER M4 ;
			RECT 0.000 135.955 80.085 136.285 ;
			LAYER M4 ;
			RECT 0.000 138.275 80.085 138.605 ;
			LAYER M4 ;
			RECT 0.000 140.595 80.085 140.925 ;
			LAYER M4 ;
			RECT 0.000 142.915 80.085 143.245 ;
			LAYER M4 ;
			RECT 0.000 145.235 80.085 145.565 ;
			LAYER M4 ;
			RECT 0.000 147.555 80.085 147.885 ;
			LAYER M4 ;
			RECT 0.000 149.905 80.085 150.210 ;
			LAYER M4 ;
			RECT 0.000 153.770 80.085 154.320 ;
			LAYER M4 ;
			RECT 0.000 154.825 80.085 155.245 ;
			LAYER M4 ;
			RECT 0.000 156.790 80.085 157.360 ;
			LAYER M4 ;
			RECT 0.000 157.490 80.085 158.060 ;
			LAYER M4 ;
			RECT 56.840 160.200 80.085 160.850 ;
			LAYER M4 ;
			RECT 0.000 161.950 80.085 162.600 ;
			LAYER M4 ;
			RECT 0.000 164.745 80.085 165.395 ;
			LAYER M4 ;
			RECT 0.000 165.545 80.085 165.855 ;
			LAYER M4 ;
			RECT 0.000 168.395 80.085 168.725 ;
			LAYER M4 ;
			RECT 0.000 170.715 80.085 171.045 ;
			LAYER M4 ;
			RECT 0.000 173.035 80.085 173.365 ;
			LAYER M4 ;
			RECT 0.000 175.355 80.085 175.685 ;
			LAYER M4 ;
			RECT 0.000 177.675 80.085 178.005 ;
			LAYER M4 ;
			RECT 0.000 179.995 80.085 180.325 ;
			LAYER M4 ;
			RECT 0.000 182.315 80.085 182.645 ;
			LAYER M4 ;
			RECT 0.000 184.635 80.085 184.965 ;
			LAYER M4 ;
			RECT 0.000 186.955 80.085 187.285 ;
			LAYER M4 ;
			RECT 0.000 189.275 80.085 189.605 ;
			LAYER M4 ;
			RECT 0.000 191.595 80.085 191.925 ;
			LAYER M4 ;
			RECT 0.000 193.915 80.085 194.245 ;
			LAYER M4 ;
			RECT 0.000 196.235 80.085 196.565 ;
			LAYER M4 ;
			RECT 0.000 198.555 80.085 198.885 ;
			LAYER M4 ;
			RECT 0.000 200.875 80.085 201.205 ;
			LAYER M4 ;
			RECT 0.000 203.195 80.085 203.525 ;
			LAYER M4 ;
			RECT 0.000 205.515 80.085 205.845 ;
			LAYER M4 ;
			RECT 0.000 207.835 80.085 208.165 ;
			LAYER M4 ;
			RECT 0.000 210.155 80.085 210.485 ;
			LAYER M4 ;
			RECT 0.000 212.475 80.085 212.805 ;
			LAYER M4 ;
			RECT 0.000 214.795 80.085 215.125 ;
			LAYER M4 ;
			RECT 0.000 217.115 80.085 217.445 ;
			LAYER M4 ;
			RECT 0.000 219.435 80.085 219.765 ;
			LAYER M4 ;
			RECT 0.000 221.755 80.085 222.085 ;
			LAYER M4 ;
			RECT 0.000 224.075 80.085 224.405 ;
			LAYER M4 ;
			RECT 0.000 226.395 80.085 226.725 ;
			LAYER M4 ;
			RECT 0.000 228.715 80.085 229.045 ;
			LAYER M4 ;
			RECT 0.000 231.035 80.085 231.365 ;
			LAYER M4 ;
			RECT 0.000 233.355 80.085 233.685 ;
			LAYER M4 ;
			RECT 0.000 235.675 80.085 236.005 ;
			LAYER M4 ;
			RECT 0.000 237.995 80.085 238.325 ;
			LAYER M4 ;
			RECT 0.000 240.315 80.085 240.645 ;
			LAYER M4 ;
			RECT 0.000 242.635 80.085 242.965 ;
			LAYER M4 ;
			RECT 0.000 244.955 80.085 245.285 ;
			LAYER M4 ;
			RECT 0.000 247.275 80.085 247.605 ;
			LAYER M4 ;
			RECT 0.000 249.595 80.085 249.925 ;
			LAYER M4 ;
			RECT 0.000 251.915 80.085 252.245 ;
			LAYER M4 ;
			RECT 0.000 254.235 80.085 254.565 ;
			LAYER M4 ;
			RECT 0.000 256.555 80.085 256.885 ;
			LAYER M4 ;
			RECT 0.000 258.875 80.085 259.205 ;
			LAYER M4 ;
			RECT 0.000 261.195 80.085 261.525 ;
			LAYER M4 ;
			RECT 0.000 263.515 80.085 263.845 ;
			LAYER M4 ;
			RECT 0.000 265.835 80.085 266.165 ;
			LAYER M4 ;
			RECT 0.000 268.155 80.085 268.485 ;
			LAYER M4 ;
			RECT 0.000 270.475 80.085 270.805 ;
			LAYER M4 ;
			RECT 0.000 272.795 80.085 273.125 ;
			LAYER M4 ;
			RECT 0.000 275.115 80.085 275.445 ;
			LAYER M4 ;
			RECT 0.000 277.435 80.085 277.765 ;
			LAYER M4 ;
			RECT 0.000 279.755 80.085 280.085 ;
			LAYER M4 ;
			RECT 0.000 282.075 80.085 282.405 ;
			LAYER M4 ;
			RECT 0.000 284.395 80.085 284.725 ;
			LAYER M4 ;
			RECT 0.000 286.715 80.085 287.045 ;
			LAYER M4 ;
			RECT 0.000 289.035 80.085 289.365 ;
			LAYER M4 ;
			RECT 0.000 291.355 80.085 291.685 ;
			LAYER M4 ;
			RECT 0.000 293.675 80.085 294.005 ;
			LAYER M4 ;
			RECT 0.000 295.995 80.085 296.325 ;
			LAYER M4 ;
			RECT 0.000 298.315 80.085 298.645 ;
			LAYER M4 ;
			RECT 0.000 300.635 80.085 300.965 ;
			LAYER M4 ;
			RECT 0.000 302.955 80.085 303.285 ;
			LAYER M4 ;
			RECT 0.000 305.275 80.085 305.605 ;
			LAYER M4 ;
			RECT 0.000 307.595 80.085 307.925 ;
			LAYER M4 ;
			RECT 0.000 309.915 80.085 310.245 ;
			LAYER M4 ;
			RECT 0.000 312.235 80.085 312.565 ;
			LAYER M4 ;
			RECT 0.000 314.555 80.085 314.885 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.000 2.805 80.085 3.185 ;
			LAYER M4 ;
			RECT 0.000 5.125 80.085 5.505 ;
			LAYER M4 ;
			RECT 0.000 7.445 80.085 7.825 ;
			LAYER M4 ;
			RECT 0.000 9.765 80.085 10.145 ;
			LAYER M4 ;
			RECT 0.000 12.085 80.085 12.465 ;
			LAYER M4 ;
			RECT 0.000 14.405 80.085 14.785 ;
			LAYER M4 ;
			RECT 0.000 16.725 80.085 17.105 ;
			LAYER M4 ;
			RECT 0.000 19.045 80.085 19.425 ;
			LAYER M4 ;
			RECT 0.000 21.365 80.085 21.745 ;
			LAYER M4 ;
			RECT 0.000 23.685 80.085 24.065 ;
			LAYER M4 ;
			RECT 0.000 26.005 80.085 26.385 ;
			LAYER M4 ;
			RECT 0.000 28.325 80.085 28.705 ;
			LAYER M4 ;
			RECT 0.000 30.645 80.085 31.025 ;
			LAYER M4 ;
			RECT 0.000 32.965 80.085 33.345 ;
			LAYER M4 ;
			RECT 0.000 35.285 80.085 35.665 ;
			LAYER M4 ;
			RECT 0.000 37.605 80.085 37.985 ;
			LAYER M4 ;
			RECT 0.000 39.925 80.085 40.305 ;
			LAYER M4 ;
			RECT 0.000 42.245 80.085 42.625 ;
			LAYER M4 ;
			RECT 0.000 44.565 80.085 44.945 ;
			LAYER M4 ;
			RECT 0.000 46.885 80.085 47.265 ;
			LAYER M4 ;
			RECT 0.000 49.205 80.085 49.585 ;
			LAYER M4 ;
			RECT 0.000 51.525 80.085 51.905 ;
			LAYER M4 ;
			RECT 0.000 53.845 80.085 54.225 ;
			LAYER M4 ;
			RECT 0.000 56.165 80.085 56.545 ;
			LAYER M4 ;
			RECT 0.000 58.485 80.085 58.865 ;
			LAYER M4 ;
			RECT 0.000 60.805 80.085 61.185 ;
			LAYER M4 ;
			RECT 0.000 63.125 80.085 63.505 ;
			LAYER M4 ;
			RECT 0.000 65.445 80.085 65.825 ;
			LAYER M4 ;
			RECT 0.000 67.765 80.085 68.145 ;
			LAYER M4 ;
			RECT 0.000 70.085 80.085 70.465 ;
			LAYER M4 ;
			RECT 0.000 72.405 80.085 72.785 ;
			LAYER M4 ;
			RECT 0.000 74.725 80.085 75.105 ;
			LAYER M4 ;
			RECT 0.000 77.045 80.085 77.425 ;
			LAYER M4 ;
			RECT 0.000 79.365 80.085 79.745 ;
			LAYER M4 ;
			RECT 0.000 81.685 80.085 82.065 ;
			LAYER M4 ;
			RECT 0.000 84.005 80.085 84.385 ;
			LAYER M4 ;
			RECT 0.000 86.325 80.085 86.705 ;
			LAYER M4 ;
			RECT 0.000 88.645 80.085 89.025 ;
			LAYER M4 ;
			RECT 0.000 90.965 80.085 91.345 ;
			LAYER M4 ;
			RECT 0.000 93.285 80.085 93.665 ;
			LAYER M4 ;
			RECT 0.000 95.605 80.085 95.985 ;
			LAYER M4 ;
			RECT 0.000 97.925 80.085 98.305 ;
			LAYER M4 ;
			RECT 0.000 100.245 80.085 100.625 ;
			LAYER M4 ;
			RECT 0.000 102.565 80.085 102.945 ;
			LAYER M4 ;
			RECT 0.000 104.885 80.085 105.265 ;
			LAYER M4 ;
			RECT 0.000 107.205 80.085 107.585 ;
			LAYER M4 ;
			RECT 0.000 109.525 80.085 109.905 ;
			LAYER M4 ;
			RECT 0.000 111.845 80.085 112.225 ;
			LAYER M4 ;
			RECT 0.000 114.165 80.085 114.545 ;
			LAYER M4 ;
			RECT 0.000 116.485 80.085 116.865 ;
			LAYER M4 ;
			RECT 0.000 118.805 80.085 119.185 ;
			LAYER M4 ;
			RECT 0.000 121.125 80.085 121.505 ;
			LAYER M4 ;
			RECT 0.000 123.445 80.085 123.825 ;
			LAYER M4 ;
			RECT 0.000 125.765 80.085 126.145 ;
			LAYER M4 ;
			RECT 0.000 128.085 80.085 128.465 ;
			LAYER M4 ;
			RECT 0.000 130.405 80.085 130.785 ;
			LAYER M4 ;
			RECT 0.000 132.725 80.085 133.105 ;
			LAYER M4 ;
			RECT 0.000 135.045 80.085 135.425 ;
			LAYER M4 ;
			RECT 0.000 137.365 80.085 137.745 ;
			LAYER M4 ;
			RECT 0.000 139.685 80.085 140.065 ;
			LAYER M4 ;
			RECT 0.000 142.005 80.085 142.385 ;
			LAYER M4 ;
			RECT 0.000 144.325 80.085 144.705 ;
			LAYER M4 ;
			RECT 0.000 146.645 80.085 147.025 ;
			LAYER M4 ;
			RECT 0.000 148.965 80.085 149.345 ;
			LAYER M4 ;
			RECT 54.215 152.230 80.085 153.010 ;
			LAYER M4 ;
			RECT 0.000 155.390 80.085 155.960 ;
			LAYER M4 ;
			RECT 0.000 156.090 80.085 156.660 ;
			LAYER M4 ;
			RECT 0.000 158.320 80.085 158.970 ;
			LAYER M4 ;
			RECT 56.840 159.400 80.085 160.050 ;
			LAYER M4 ;
			RECT 0.000 161.230 80.085 161.800 ;
			LAYER M4 ;
			RECT 0.000 169.805 80.085 170.185 ;
			LAYER M4 ;
			RECT 0.000 172.125 80.085 172.505 ;
			LAYER M4 ;
			RECT 0.000 174.445 80.085 174.825 ;
			LAYER M4 ;
			RECT 0.000 176.765 80.085 177.145 ;
			LAYER M4 ;
			RECT 0.000 179.085 80.085 179.465 ;
			LAYER M4 ;
			RECT 0.000 181.405 80.085 181.785 ;
			LAYER M4 ;
			RECT 0.000 183.725 80.085 184.105 ;
			LAYER M4 ;
			RECT 0.000 186.045 80.085 186.425 ;
			LAYER M4 ;
			RECT 0.000 188.365 80.085 188.745 ;
			LAYER M4 ;
			RECT 0.000 190.685 80.085 191.065 ;
			LAYER M4 ;
			RECT 0.000 193.005 80.085 193.385 ;
			LAYER M4 ;
			RECT 0.000 195.325 80.085 195.705 ;
			LAYER M4 ;
			RECT 0.000 197.645 80.085 198.025 ;
			LAYER M4 ;
			RECT 0.000 199.965 80.085 200.345 ;
			LAYER M4 ;
			RECT 0.000 202.285 80.085 202.665 ;
			LAYER M4 ;
			RECT 0.000 204.605 80.085 204.985 ;
			LAYER M4 ;
			RECT 0.000 206.925 80.085 207.305 ;
			LAYER M4 ;
			RECT 0.000 209.245 80.085 209.625 ;
			LAYER M4 ;
			RECT 0.000 211.565 80.085 211.945 ;
			LAYER M4 ;
			RECT 0.000 213.885 80.085 214.265 ;
			LAYER M4 ;
			RECT 0.000 216.205 80.085 216.585 ;
			LAYER M4 ;
			RECT 0.000 218.525 80.085 218.905 ;
			LAYER M4 ;
			RECT 0.000 220.845 80.085 221.225 ;
			LAYER M4 ;
			RECT 0.000 223.165 80.085 223.545 ;
			LAYER M4 ;
			RECT 0.000 225.485 80.085 225.865 ;
			LAYER M4 ;
			RECT 0.000 227.805 80.085 228.185 ;
			LAYER M4 ;
			RECT 0.000 230.125 80.085 230.505 ;
			LAYER M4 ;
			RECT 0.000 232.445 80.085 232.825 ;
			LAYER M4 ;
			RECT 0.000 234.765 80.085 235.145 ;
			LAYER M4 ;
			RECT 0.000 237.085 80.085 237.465 ;
			LAYER M4 ;
			RECT 0.000 239.405 80.085 239.785 ;
			LAYER M4 ;
			RECT 0.000 241.725 80.085 242.105 ;
			LAYER M4 ;
			RECT 0.000 244.045 80.085 244.425 ;
			LAYER M4 ;
			RECT 0.000 246.365 80.085 246.745 ;
			LAYER M4 ;
			RECT 0.000 248.685 80.085 249.065 ;
			LAYER M4 ;
			RECT 0.000 251.005 80.085 251.385 ;
			LAYER M4 ;
			RECT 0.000 253.325 80.085 253.705 ;
			LAYER M4 ;
			RECT 0.000 255.645 80.085 256.025 ;
			LAYER M4 ;
			RECT 0.000 257.965 80.085 258.345 ;
			LAYER M4 ;
			RECT 0.000 260.285 80.085 260.665 ;
			LAYER M4 ;
			RECT 0.000 262.605 80.085 262.985 ;
			LAYER M4 ;
			RECT 0.000 264.925 80.085 265.305 ;
			LAYER M4 ;
			RECT 0.000 267.245 80.085 267.625 ;
			LAYER M4 ;
			RECT 0.000 269.565 80.085 269.945 ;
			LAYER M4 ;
			RECT 0.000 271.885 80.085 272.265 ;
			LAYER M4 ;
			RECT 0.000 274.205 80.085 274.585 ;
			LAYER M4 ;
			RECT 0.000 276.525 80.085 276.905 ;
			LAYER M4 ;
			RECT 0.000 278.845 80.085 279.225 ;
			LAYER M4 ;
			RECT 0.000 281.165 80.085 281.545 ;
			LAYER M4 ;
			RECT 0.000 283.485 80.085 283.865 ;
			LAYER M4 ;
			RECT 0.000 285.805 80.085 286.185 ;
			LAYER M4 ;
			RECT 0.000 288.125 80.085 288.505 ;
			LAYER M4 ;
			RECT 0.000 290.445 80.085 290.825 ;
			LAYER M4 ;
			RECT 0.000 292.765 80.085 293.145 ;
			LAYER M4 ;
			RECT 0.000 295.085 80.085 295.465 ;
			LAYER M4 ;
			RECT 0.000 297.405 80.085 297.785 ;
			LAYER M4 ;
			RECT 0.000 299.725 80.085 300.105 ;
			LAYER M4 ;
			RECT 0.000 302.045 80.085 302.425 ;
			LAYER M4 ;
			RECT 0.000 304.365 80.085 304.745 ;
			LAYER M4 ;
			RECT 0.000 306.685 80.085 307.065 ;
			LAYER M4 ;
			RECT 0.000 309.005 80.085 309.385 ;
			LAYER M4 ;
			RECT 0.000 311.325 80.085 311.705 ;
			LAYER M4 ;
			RECT 0.000 313.645 80.085 314.025 ;
			LAYER M4 ;
			RECT 0.000 315.965 80.085 316.345 ;
		END
	END VSS

	PIN WEBA
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 162.365 80.475 162.515 ;
			LAYER M1 ;
			RECT 80.295 162.365 80.475 162.515 ;
			LAYER M3 ;
			RECT 80.295 162.365 80.475 162.515 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.170000 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.166700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.530800 LAYER M2 ;
		ANTENNAMAXAREACAR 15.783300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.122900 LAYER M3 ;
		ANTENNAMAXAREACAR 17.051300 LAYER M3 ;
	END WEBA

	PIN WEBB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.295 162.695 80.475 162.845 ;
			LAYER M1 ;
			RECT 80.295 162.695 80.475 162.845 ;
			LAYER M2 ;
			RECT 80.295 162.695 80.475 162.845 ;
		END
		ANTENNAGATEAREA 0.022500 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.088700 LAYER M1 ;
		ANTENNAMAXAREACAR 1.788900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.288900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.022500 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.465500 LAYER M2 ;
		ANTENNAMAXAREACAR 20.633300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.577800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.022500 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.080200 LAYER M3 ;
		ANTENNAMAXAREACAR 21.833300 LAYER M3 ;
	END WEBB

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 167.275 80.475 167.425 ;
			LAYER M3 ;
			RECT 80.295 167.275 80.475 167.425 ;
			LAYER M1 ;
			RECT 80.295 167.275 80.475 167.425 ;
		END
		ANTENNAGATEAREA 0.022500 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.073500 LAYER M1 ;
		ANTENNAMAXAREACAR 1.111100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.288900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.022500 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.383200 LAYER M2 ;
		ANTENNAMAXAREACAR 17.766700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.577800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.022500 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.202700 LAYER M3 ;
		ANTENNAMAXAREACAR 18.966700 LAYER M3 ;
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.295 166.290 80.475 166.440 ;
			LAYER M3 ;
			RECT 80.295 166.290 80.475 166.440 ;
			LAYER M1 ;
			RECT 80.295 166.290 80.475 166.440 ;
		END
		ANTENNAGATEAREA 0.022500 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.073500 LAYER M1 ;
		ANTENNAMAXAREACAR 1.111100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.288900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.022500 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.383200 LAYER M2 ;
		ANTENNAMAXAREACAR 17.766700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.577800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.022500 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.202700 LAYER M3 ;
		ANTENNAMAXAREACAR 18.966700 LAYER M3 ;
	END WTSEL[1]

	OBS
		# Promoted blockages
		LAYER M2 ;
		RECT 80.295 316.575 80.475 317.690 ;
		LAYER VIA3 ;
		RECT 80.295 315.915 80.475 315.935 ;
		LAYER M1 ;
		RECT 80.295 315.230 80.475 315.625 ;
		LAYER VIA3 ;
		RECT 80.295 315.250 80.475 315.605 ;
		LAYER M2 ;
		RECT 80.295 266.530 80.475 266.885 ;
		LAYER M3 ;
		RECT 80.295 266.530 80.475 266.885 ;
		LAYER M2 ;
		RECT 80.295 265.535 80.475 266.220 ;
		LAYER M3 ;
		RECT 80.295 265.535 80.475 266.220 ;
		LAYER VIA3 ;
		RECT 80.295 266.530 80.475 266.885 ;
		LAYER M2 ;
		RECT 80.295 267.195 80.475 267.215 ;
		LAYER M2 ;
		RECT 80.295 267.525 80.475 267.545 ;
		LAYER M2 ;
		RECT 80.295 267.855 80.475 268.540 ;
		LAYER M3 ;
		RECT 80.295 267.855 80.475 268.540 ;
		LAYER M3 ;
		RECT 80.295 267.525 80.475 267.545 ;
		LAYER M3 ;
		RECT 80.295 267.195 80.475 267.215 ;
		LAYER VIA3 ;
		RECT 80.295 267.195 80.475 267.215 ;
		LAYER M1 ;
		RECT 80.295 267.835 80.475 268.560 ;
		LAYER VIA3 ;
		RECT 80.295 309.615 80.475 310.300 ;
		LAYER M1 ;
		RECT 80.295 309.595 80.475 310.320 ;
		LAYER M2 ;
		RECT 80.295 309.285 80.475 309.305 ;
		LAYER VIA3 ;
		RECT 80.295 311.935 80.475 312.620 ;
		LAYER M1 ;
		RECT 80.295 311.915 80.475 312.640 ;
		LAYER VIA3 ;
		RECT 80.295 302.655 80.475 303.340 ;
		LAYER VIA3 ;
		RECT 80.295 303.650 80.475 304.005 ;
		LAYER M3 ;
		RECT 80.295 299.675 80.475 299.695 ;
		LAYER VIA3 ;
		RECT 80.295 299.675 80.475 299.695 ;
		LAYER M1 ;
		RECT 80.295 301.310 80.475 301.705 ;
		LAYER M2 ;
		RECT 80.295 295.035 80.475 295.055 ;
		LAYER M2 ;
		RECT 80.295 294.370 80.475 294.725 ;
		LAYER M3 ;
		RECT 80.295 294.370 80.475 294.725 ;
		LAYER M1 ;
		RECT 80.295 294.350 80.475 294.745 ;
		LAYER M3 ;
		RECT 80.295 295.035 80.475 295.055 ;
		LAYER VIA3 ;
		RECT 80.295 294.370 80.475 294.725 ;
		LAYER VIA3 ;
		RECT 80.295 297.685 80.475 297.705 ;
		LAYER M2 ;
		RECT 80.295 293.375 80.475 294.060 ;
		LAYER M3 ;
		RECT 80.295 293.375 80.475 294.060 ;
		LAYER M1 ;
		RECT 80.295 281.425 80.475 281.485 ;
		LAYER M1 ;
		RECT 80.295 281.095 80.475 281.155 ;
		LAYER M1 ;
		RECT 80.295 280.430 80.475 280.825 ;
		LAYER M2 ;
		RECT 80.295 285.090 80.475 285.445 ;
		LAYER M2 ;
		RECT 80.295 293.045 80.475 293.065 ;
		LAYER M1 ;
		RECT 80.295 293.025 80.475 293.085 ;
		LAYER M3 ;
		RECT 80.295 292.715 80.475 292.735 ;
		LAYER M1 ;
		RECT 80.295 292.695 80.475 292.755 ;
		LAYER M1 ;
		RECT 80.295 292.030 80.475 292.425 ;
		LAYER VIA3 ;
		RECT 80.295 291.055 80.475 291.740 ;
		LAYER M1 ;
		RECT 80.295 0.000 80.475 1.800 ;
		LAYER M1 ;
		RECT 80.295 2.735 80.475 2.795 ;
		LAYER M2 ;
		RECT 80.295 2.755 80.475 2.775 ;
		LAYER M3 ;
		RECT 80.295 2.755 80.475 2.775 ;
		LAYER VIA3 ;
		RECT 80.295 2.755 80.475 2.775 ;
		LAYER M1 ;
		RECT 80.295 3.065 80.475 3.125 ;
		LAYER M2 ;
		RECT 80.295 0.000 80.475 1.780 ;
		LAYER M3 ;
		RECT 80.295 0.000 80.475 1.780 ;
		LAYER VIA3 ;
		RECT 80.295 0.000 80.475 1.780 ;
		LAYER M1 ;
		RECT 80.295 9.695 80.475 9.755 ;
		LAYER M2 ;
		RECT 80.295 10.045 80.475 10.065 ;
		LAYER M2 ;
		RECT 80.295 10.375 80.475 11.060 ;
		LAYER M2 ;
		RECT 80.295 11.370 80.475 11.725 ;
		LAYER M2 ;
		RECT 80.295 2.090 80.475 2.445 ;
		LAYER M3 ;
		RECT 80.295 2.090 80.475 2.445 ;
		LAYER VIA3 ;
		RECT 80.295 2.090 80.475 2.445 ;
		LAYER M1 ;
		RECT 80.295 2.070 80.475 2.465 ;
		LAYER M1 ;
		RECT 80.295 237.345 80.475 237.405 ;
		LAYER VIA3 ;
		RECT 80.295 237.035 80.475 237.055 ;
		LAYER M2 ;
		RECT 80.295 237.035 80.475 237.055 ;
		LAYER M3 ;
		RECT 80.295 237.035 80.475 237.055 ;
		LAYER VIA3 ;
		RECT 80.295 236.370 80.475 236.725 ;
		LAYER VIA3 ;
		RECT 80.295 235.375 80.475 236.060 ;
		LAYER VIA3 ;
		RECT 80.295 235.045 80.475 235.065 ;
		LAYER M3 ;
		RECT 80.295 236.370 80.475 236.725 ;
		LAYER M3 ;
		RECT 80.295 235.375 80.475 236.060 ;
		LAYER M3 ;
		RECT 80.295 233.055 80.475 233.740 ;
		LAYER M3 ;
		RECT 80.295 234.715 80.475 234.735 ;
		LAYER M3 ;
		RECT 80.295 234.050 80.475 234.405 ;
		LAYER M2 ;
		RECT 80.295 237.365 80.475 237.385 ;
		LAYER M2 ;
		RECT 80.295 239.355 80.475 239.375 ;
		LAYER M3 ;
		RECT 80.295 239.355 80.475 239.375 ;
		LAYER M1 ;
		RECT 80.295 237.675 80.475 238.400 ;
		LAYER M2 ;
		RECT 80.295 239.685 80.475 239.705 ;
		LAYER M1 ;
		RECT 80.295 239.665 80.475 239.725 ;
		LAYER M1 ;
		RECT 80.295 239.335 80.475 239.395 ;
		LAYER M2 ;
		RECT 80.295 240.015 80.475 240.700 ;
		LAYER M3 ;
		RECT 80.295 239.685 80.475 239.705 ;
		LAYER M1 ;
		RECT 80.295 240.990 80.475 241.385 ;
		LAYER M2 ;
		RECT 80.295 241.675 80.475 241.695 ;
		LAYER M2 ;
		RECT 80.295 244.325 80.475 244.345 ;
		LAYER VIA3 ;
		RECT 80.295 243.995 80.475 244.015 ;
		LAYER VIA3 ;
		RECT 80.295 243.330 80.475 243.685 ;
		LAYER VIA3 ;
		RECT 80.295 242.335 80.475 243.020 ;
		LAYER M3 ;
		RECT 80.295 244.325 80.475 244.345 ;
		LAYER VIA3 ;
		RECT 80.295 244.325 80.475 244.345 ;
		LAYER VIA3 ;
		RECT 80.295 242.005 80.475 242.025 ;
		LAYER M3 ;
		RECT 80.295 240.015 80.475 240.700 ;
		LAYER M1 ;
		RECT 80.295 239.995 80.475 240.720 ;
		LAYER M2 ;
		RECT 80.295 241.010 80.475 241.365 ;
		LAYER M3 ;
		RECT 80.295 241.010 80.475 241.365 ;
		LAYER M1 ;
		RECT 80.295 225.745 80.475 225.805 ;
		LAYER M3 ;
		RECT 80.295 219.135 80.475 219.820 ;
		LAYER M1 ;
		RECT 80.295 220.110 80.475 220.505 ;
		LAYER M3 ;
		RECT 80.295 170.120 80.475 170.800 ;
		LAYER M1 ;
		RECT 80.295 170.100 80.475 170.820 ;
		LAYER VIA3 ;
		RECT 80.295 169.160 80.475 169.810 ;
		LAYER M1 ;
		RECT 80.295 169.140 80.475 169.830 ;
		LAYER M2 ;
		RECT 80.295 163.585 80.475 163.900 ;
		LAYER M3 ;
		RECT 80.295 163.585 80.475 163.900 ;
		LAYER M1 ;
		RECT 80.295 163.565 80.475 163.920 ;
		LAYER M2 ;
		RECT 80.295 163.255 80.475 163.275 ;
		LAYER M2 ;
		RECT 80.295 201.570 80.475 201.925 ;
		LAYER M1 ;
		RECT 80.295 202.215 80.475 202.275 ;
		LAYER M1 ;
		RECT 80.295 168.810 80.475 168.870 ;
		LAYER M3 ;
		RECT 80.295 225.435 80.475 225.455 ;
		LAYER VIA3 ;
		RECT 80.295 220.130 80.475 220.485 ;
		LAYER M2 ;
		RECT 80.295 220.130 80.475 220.485 ;
		LAYER M1 ;
		RECT 80.295 222.430 80.475 222.825 ;
		LAYER M2 ;
		RECT 80.295 222.450 80.475 222.805 ;
		LAYER M1 ;
		RECT 80.295 225.415 80.475 225.475 ;
		LAYER M3 ;
		RECT 80.295 223.775 80.475 224.460 ;
		LAYER M2 ;
		RECT 80.295 223.445 80.475 223.465 ;
		LAYER M2 ;
		RECT 80.295 223.115 80.475 223.135 ;
		LAYER M2 ;
		RECT 80.295 168.500 80.475 168.520 ;
		LAYER VIA3 ;
		RECT 80.295 168.500 80.475 168.520 ;
		LAYER VIA3 ;
		RECT 80.295 167.505 80.475 168.190 ;
		LAYER M2 ;
		RECT 80.295 167.505 80.475 168.190 ;
		LAYER M3 ;
		RECT 80.295 167.505 80.475 168.190 ;
		LAYER M2 ;
		RECT 80.295 166.520 80.475 166.540 ;
		LAYER M2 ;
		RECT 80.295 164.870 80.475 166.210 ;
		LAYER VIA3 ;
		RECT 80.295 164.540 80.475 164.560 ;
		LAYER VIA3 ;
		RECT 80.295 164.210 80.475 164.230 ;
		LAYER VIA3 ;
		RECT 80.295 166.520 80.475 166.540 ;
		LAYER VIA3 ;
		RECT 80.295 168.830 80.475 168.850 ;
		LAYER M2 ;
		RECT 80.295 168.830 80.475 168.850 ;
		LAYER M1 ;
		RECT 80.295 168.480 80.475 168.540 ;
		LAYER M1 ;
		RECT 80.295 167.485 80.475 168.210 ;
		LAYER M3 ;
		RECT 80.295 168.830 80.475 168.850 ;
		LAYER M3 ;
		RECT 80.295 168.500 80.475 168.520 ;
		LAYER VIA3 ;
		RECT 80.295 163.255 80.475 163.275 ;
		LAYER M3 ;
		RECT 80.295 163.255 80.475 163.275 ;
		LAYER M1 ;
		RECT 80.295 167.160 80.475 167.215 ;
		LAYER VIA3 ;
		RECT 80.295 163.585 80.475 163.900 ;
		LAYER M1 ;
		RECT 80.295 164.190 80.475 164.250 ;
		LAYER M1 ;
		RECT 80.295 166.830 80.475 166.890 ;
		LAYER M1 ;
		RECT 80.295 166.500 80.475 166.560 ;
		LAYER VIA3 ;
		RECT 80.295 167.180 80.475 167.195 ;
		LAYER M2 ;
		RECT 80.295 167.180 80.475 167.195 ;
		LAYER M3 ;
		RECT 80.295 167.180 80.475 167.195 ;
		LAYER M1 ;
		RECT 80.295 232.705 80.475 232.765 ;
		LAYER M2 ;
		RECT 80.295 232.725 80.475 232.745 ;
		LAYER M2 ;
		RECT 80.295 230.405 80.475 230.425 ;
		LAYER M3 ;
		RECT 80.295 232.725 80.475 232.745 ;
		LAYER M1 ;
		RECT 80.295 232.375 80.475 232.435 ;
		LAYER M2 ;
		RECT 80.295 232.395 80.475 232.415 ;
		LAYER M2 ;
		RECT 80.295 231.730 80.475 232.085 ;
		LAYER M2 ;
		RECT 80.295 230.735 80.475 231.420 ;
		LAYER VIA3 ;
		RECT 80.295 232.395 80.475 232.415 ;
		LAYER VIA3 ;
		RECT 80.295 230.735 80.475 231.420 ;
		LAYER M1 ;
		RECT 80.295 230.385 80.475 230.445 ;
		LAYER VIA3 ;
		RECT 80.295 230.405 80.475 230.425 ;
		LAYER M1 ;
		RECT 80.295 229.390 80.475 229.785 ;
		LAYER M2 ;
		RECT 80.295 228.415 80.475 229.100 ;
		LAYER VIA3 ;
		RECT 80.295 228.415 80.475 229.100 ;
		LAYER VIA3 ;
		RECT 80.295 228.085 80.475 228.105 ;
		LAYER VIA3 ;
		RECT 80.295 227.755 80.475 227.775 ;
		LAYER VIA3 ;
		RECT 80.295 227.090 80.475 227.445 ;
		LAYER M3 ;
		RECT 80.295 227.090 80.475 227.445 ;
		LAYER M2 ;
		RECT 80.295 230.075 80.475 230.095 ;
		LAYER VIA3 ;
		RECT 80.295 230.075 80.475 230.095 ;
		LAYER M1 ;
		RECT 80.295 230.055 80.475 230.115 ;
		LAYER VIA3 ;
		RECT 80.295 229.410 80.475 229.765 ;
		LAYER M2 ;
		RECT 80.295 237.695 80.475 238.380 ;
		LAYER M2 ;
		RECT 80.295 238.690 80.475 239.045 ;
		LAYER M1 ;
		RECT 80.295 238.670 80.475 239.065 ;
		LAYER M2 ;
		RECT 80.295 245.650 80.475 246.005 ;
		LAYER VIA3 ;
		RECT 80.295 245.650 80.475 246.005 ;
		LAYER M3 ;
		RECT 80.295 242.335 80.475 243.020 ;
		LAYER M3 ;
		RECT 80.295 245.650 80.475 246.005 ;
		LAYER M2 ;
		RECT 80.295 242.335 80.475 243.020 ;
		LAYER M2 ;
		RECT 80.295 242.005 80.475 242.025 ;
		LAYER M3 ;
		RECT 80.295 242.005 80.475 242.025 ;
		LAYER M3 ;
		RECT 80.295 17.005 80.475 17.025 ;
		LAYER M2 ;
		RECT 80.295 17.005 80.475 17.025 ;
		LAYER VIA3 ;
		RECT 80.295 26.615 80.475 27.300 ;
		LAYER M3 ;
		RECT 80.295 29.930 80.475 30.285 ;
		LAYER VIA3 ;
		RECT 80.295 29.930 80.475 30.285 ;
		LAYER M3 ;
		RECT 80.295 28.935 80.475 29.620 ;
		LAYER VIA3 ;
		RECT 80.295 28.935 80.475 29.620 ;
		LAYER M2 ;
		RECT 80.295 29.930 80.475 30.285 ;
		LAYER M1 ;
		RECT 80.295 31.235 80.475 31.960 ;
		LAYER VIA3 ;
		RECT 80.295 31.255 80.475 31.940 ;
		LAYER M2 ;
		RECT 80.295 30.595 80.475 30.615 ;
		LAYER M3 ;
		RECT 80.295 30.595 80.475 30.615 ;
		LAYER M2 ;
		RECT 80.295 31.255 80.475 31.940 ;
		LAYER M2 ;
		RECT 80.295 63.075 80.475 63.095 ;
		LAYER M2 ;
		RECT 80.295 27.610 80.475 27.965 ;
		LAYER VIA3 ;
		RECT 80.295 27.610 80.475 27.965 ;
		LAYER M3 ;
		RECT 80.295 28.605 80.475 28.625 ;
		LAYER VIA3 ;
		RECT 80.295 28.605 80.475 28.625 ;
		LAYER M1 ;
		RECT 80.295 18.310 80.475 18.705 ;
		LAYER M2 ;
		RECT 80.295 18.995 80.475 19.015 ;
		LAYER M3 ;
		RECT 80.295 26.285 80.475 26.305 ;
		LAYER M2 ;
		RECT 80.295 26.615 80.475 27.300 ;
		LAYER M3 ;
		RECT 80.295 38.215 80.475 38.900 ;
		LAYER M1 ;
		RECT 80.295 32.230 80.475 32.625 ;
		LAYER M3 ;
		RECT 80.295 32.250 80.475 32.605 ;
		LAYER M1 ;
		RECT 80.295 114.755 80.475 115.480 ;
		LAYER VIA3 ;
		RECT 80.295 114.775 80.475 115.460 ;
		LAYER VIA3 ;
		RECT 80.295 100.525 80.475 100.545 ;
		LAYER VIA3 ;
		RECT 80.295 98.535 80.475 99.220 ;
		LAYER M2 ;
		RECT 80.295 114.775 80.475 115.460 ;
		LAYER VIA3 ;
		RECT 80.295 102.515 80.475 102.535 ;
		LAYER VIA3 ;
		RECT 80.295 101.850 80.475 102.205 ;
		LAYER VIA3 ;
		RECT 80.295 100.855 80.475 101.540 ;
		LAYER VIA3 ;
		RECT 80.295 114.445 80.475 114.465 ;
		LAYER M1 ;
		RECT 80.295 112.435 80.475 113.160 ;
		LAYER M2 ;
		RECT 80.295 112.125 80.475 112.145 ;
		LAYER M1 ;
		RECT 80.295 112.105 80.475 112.165 ;
		LAYER M1 ;
		RECT 80.295 114.095 80.475 114.155 ;
		LAYER M3 ;
		RECT 80.295 114.445 80.475 114.465 ;
		LAYER M2 ;
		RECT 80.295 111.795 80.475 111.815 ;
		LAYER M1 ;
		RECT 80.295 111.775 80.475 111.835 ;
		LAYER VIA3 ;
		RECT 80.295 111.795 80.475 111.815 ;
		LAYER M1 ;
		RECT 80.295 115.750 80.475 116.145 ;
		LAYER M2 ;
		RECT 80.295 115.770 80.475 116.125 ;
		LAYER M3 ;
		RECT 80.295 115.770 80.475 116.125 ;
		LAYER M2 ;
		RECT 80.295 109.475 80.475 109.495 ;
		LAYER M1 ;
		RECT 80.295 110.115 80.475 110.840 ;
		LAYER VIA3 ;
		RECT 80.295 110.135 80.475 110.820 ;
		LAYER M1 ;
		RECT 80.295 311.585 80.475 311.645 ;
		LAYER M2 ;
		RECT 80.295 311.605 80.475 311.625 ;
		LAYER M3 ;
		RECT 80.295 311.605 80.475 311.625 ;
		LAYER VIA3 ;
		RECT 80.295 311.275 80.475 311.295 ;
		LAYER M2 ;
		RECT 80.295 304.975 80.475 305.660 ;
		LAYER VIA3 ;
		RECT 80.295 304.975 80.475 305.660 ;
		LAYER M1 ;
		RECT 80.295 296.670 80.475 297.065 ;
		LAYER M3 ;
		RECT 80.295 295.695 80.475 296.380 ;
		LAYER VIA3 ;
		RECT 80.295 295.695 80.475 296.380 ;
		LAYER M1 ;
		RECT 80.295 295.675 80.475 296.400 ;
		LAYER M2 ;
		RECT 80.295 297.355 80.475 297.375 ;
		LAYER M3 ;
		RECT 80.295 297.355 80.475 297.375 ;
		LAYER VIA3 ;
		RECT 80.295 297.355 80.475 297.375 ;
		LAYER M2 ;
		RECT 80.295 296.690 80.475 297.045 ;
		LAYER M3 ;
		RECT 80.295 296.690 80.475 297.045 ;
		LAYER VIA3 ;
		RECT 80.295 296.690 80.475 297.045 ;
		LAYER M3 ;
		RECT 80.295 272.495 80.475 273.180 ;
		LAYER M2 ;
		RECT 80.295 273.490 80.475 273.845 ;
		LAYER VIA3 ;
		RECT 80.295 273.490 80.475 273.845 ;
		LAYER M1 ;
		RECT 80.295 273.470 80.475 273.865 ;
		LAYER M1 ;
		RECT 80.295 287.390 80.475 287.785 ;
		LAYER VIA3 ;
		RECT 80.295 285.090 80.475 285.445 ;
		LAYER M1 ;
		RECT 80.295 285.070 80.475 285.465 ;
		LAYER VIA3 ;
		RECT 80.295 290.725 80.475 290.745 ;
		LAYER M3 ;
		RECT 80.295 290.725 80.475 290.745 ;
		LAYER M1 ;
		RECT 80.295 291.035 80.475 291.760 ;
		LAYER VIA3 ;
		RECT 80.295 292.715 80.475 292.735 ;
		LAYER M3 ;
		RECT 80.295 288.405 80.475 288.425 ;
		LAYER M3 ;
		RECT 80.295 288.735 80.475 289.420 ;
		LAYER VIA3 ;
		RECT 80.295 293.375 80.475 294.060 ;
		LAYER M1 ;
		RECT 80.295 293.355 80.475 294.080 ;
		LAYER VIA3 ;
		RECT 80.295 306.965 80.475 306.985 ;
		LAYER M3 ;
		RECT 80.295 306.965 80.475 306.985 ;
		LAYER M3 ;
		RECT 80.295 309.285 80.475 309.305 ;
		LAYER M2 ;
		RECT 80.295 305.970 80.475 306.325 ;
		LAYER M3 ;
		RECT 80.295 305.970 80.475 306.325 ;
		LAYER VIA3 ;
		RECT 80.295 305.970 80.475 306.325 ;
		LAYER M1 ;
		RECT 80.295 305.950 80.475 306.345 ;
		LAYER VIA3 ;
		RECT 80.295 301.995 80.475 302.015 ;
		LAYER VIA3 ;
		RECT 80.295 301.330 80.475 301.685 ;
		LAYER VIA3 ;
		RECT 80.295 298.015 80.475 298.700 ;
		LAYER M1 ;
		RECT 80.295 297.995 80.475 298.720 ;
		LAYER VIA3 ;
		RECT 80.295 304.645 80.475 304.665 ;
		LAYER M2 ;
		RECT 80.295 297.685 80.475 297.705 ;
		LAYER M3 ;
		RECT 80.295 297.685 80.475 297.705 ;
		LAYER M3 ;
		RECT 80.295 272.165 80.475 272.185 ;
		LAYER M2 ;
		RECT 80.295 274.155 80.475 274.175 ;
		LAYER M3 ;
		RECT 80.295 274.155 80.475 274.175 ;
		LAYER M2 ;
		RECT 80.295 274.485 80.475 274.505 ;
		LAYER VIA3 ;
		RECT 80.295 274.155 80.475 274.175 ;
		LAYER M3 ;
		RECT 80.295 274.485 80.475 274.505 ;
		LAYER VIA3 ;
		RECT 80.295 272.165 80.475 272.185 ;
		LAYER M3 ;
		RECT 80.295 278.130 80.475 278.485 ;
		LAYER VIA3 ;
		RECT 80.295 278.130 80.475 278.485 ;
		LAYER VIA3 ;
		RECT 80.295 281.775 80.475 282.460 ;
		LAYER M1 ;
		RECT 80.295 281.755 80.475 282.480 ;
		LAYER VIA3 ;
		RECT 80.295 282.770 80.475 283.125 ;
		LAYER M1 ;
		RECT 80.295 282.750 80.475 283.145 ;
		LAYER M2 ;
		RECT 80.295 282.770 80.475 283.125 ;
		LAYER M3 ;
		RECT 80.295 282.770 80.475 283.125 ;
		LAYER M3 ;
		RECT 80.295 281.115 80.475 281.135 ;
		LAYER M3 ;
		RECT 80.295 284.095 80.475 284.780 ;
		LAYER M1 ;
		RECT 80.295 284.075 80.475 284.800 ;
		LAYER VIA3 ;
		RECT 80.295 281.115 80.475 281.135 ;
		LAYER VIA3 ;
		RECT 80.295 281.445 80.475 281.465 ;
		LAYER M1 ;
		RECT 80.295 274.795 80.475 275.520 ;
		LAYER M3 ;
		RECT 80.295 277.135 80.475 277.820 ;
		LAYER M2 ;
		RECT 80.295 277.135 80.475 277.820 ;
		LAYER VIA3 ;
		RECT 80.295 274.815 80.475 275.500 ;
		LAYER VIA3 ;
		RECT 80.295 277.135 80.475 277.820 ;
		LAYER VIA3 ;
		RECT 80.295 275.810 80.475 276.165 ;
		LAYER M1 ;
		RECT 80.295 275.790 80.475 276.185 ;
		LAYER M3 ;
		RECT 80.295 276.475 80.475 276.495 ;
		LAYER VIA3 ;
		RECT 80.295 276.475 80.475 276.495 ;
		LAYER M1 ;
		RECT 80.295 311.255 80.475 311.315 ;
		LAYER M2 ;
		RECT 80.295 308.290 80.475 308.645 ;
		LAYER M3 ;
		RECT 80.295 308.290 80.475 308.645 ;
		LAYER M1 ;
		RECT 80.295 308.270 80.475 308.665 ;
		LAYER M2 ;
		RECT 80.295 252.610 80.475 252.965 ;
		LAYER M1 ;
		RECT 80.295 252.590 80.475 252.985 ;
		LAYER M2 ;
		RECT 80.295 253.275 80.475 253.295 ;
		LAYER M3 ;
		RECT 80.295 253.275 80.475 253.295 ;
		LAYER M3 ;
		RECT 80.295 252.610 80.475 252.965 ;
		LAYER M1 ;
		RECT 80.295 251.265 80.475 251.325 ;
		LAYER M2 ;
		RECT 80.295 251.285 80.475 251.305 ;
		LAYER M2 ;
		RECT 80.295 250.955 80.475 250.975 ;
		LAYER M1 ;
		RECT 80.295 250.935 80.475 250.995 ;
		LAYER M3 ;
		RECT 80.295 258.575 80.475 259.260 ;
		LAYER M1 ;
		RECT 80.295 260.875 80.475 261.600 ;
		LAYER M1 ;
		RECT 80.295 283.415 80.475 283.475 ;
		LAYER M3 ;
		RECT 80.295 271.835 80.475 271.855 ;
		LAYER M3 ;
		RECT 80.295 260.895 80.475 261.580 ;
		LAYER M2 ;
		RECT 80.295 268.850 80.475 269.205 ;
		LAYER M3 ;
		RECT 80.295 268.850 80.475 269.205 ;
		LAYER M1 ;
		RECT 80.295 269.495 80.475 269.555 ;
		LAYER M1 ;
		RECT 80.295 268.830 80.475 269.225 ;
		LAYER M3 ;
		RECT 80.295 279.455 80.475 280.140 ;
		LAYER VIA3 ;
		RECT 80.295 274.485 80.475 274.505 ;
		LAYER M3 ;
		RECT 80.295 273.490 80.475 273.845 ;
		LAYER M1 ;
		RECT 80.295 279.435 80.475 280.160 ;
		LAYER M3 ;
		RECT 80.295 283.435 80.475 283.455 ;
		LAYER VIA3 ;
		RECT 80.295 283.435 80.475 283.455 ;
		LAYER VIA3 ;
		RECT 80.295 279.455 80.475 280.140 ;
		LAYER M2 ;
		RECT 80.295 269.845 80.475 269.865 ;
		LAYER VIA3 ;
		RECT 80.295 271.835 80.475 271.855 ;
		LAYER M3 ;
		RECT 80.295 271.170 80.475 271.525 ;
		LAYER VIA3 ;
		RECT 80.295 271.170 80.475 271.525 ;
		LAYER M1 ;
		RECT 80.295 271.150 80.475 271.545 ;
		LAYER VIA3 ;
		RECT 80.295 310.610 80.475 310.965 ;
		LAYER M1 ;
		RECT 80.295 290.375 80.475 290.435 ;
		LAYER VIA3 ;
		RECT 80.295 290.395 80.475 290.415 ;
		LAYER VIA3 ;
		RECT 80.295 309.285 80.475 309.305 ;
		LAYER M1 ;
		RECT 80.295 290.705 80.475 290.765 ;
		LAYER M2 ;
		RECT 80.295 295.695 80.475 296.380 ;
		LAYER VIA3 ;
		RECT 80.295 293.045 80.475 293.065 ;
		LAYER M3 ;
		RECT 80.295 293.045 80.475 293.065 ;
		LAYER M2 ;
		RECT 80.295 295.365 80.475 295.385 ;
		LAYER M3 ;
		RECT 80.295 295.365 80.475 295.385 ;
		LAYER VIA3 ;
		RECT 80.295 295.365 80.475 295.385 ;
		LAYER VIA3 ;
		RECT 80.295 295.035 80.475 295.055 ;
		LAYER M1 ;
		RECT 80.295 286.395 80.475 287.120 ;
		LAYER VIA3 ;
		RECT 80.295 286.085 80.475 286.105 ;
		LAYER VIA3 ;
		RECT 80.295 287.410 80.475 287.765 ;
		LAYER VIA3 ;
		RECT 80.295 288.075 80.475 288.095 ;
		LAYER M3 ;
		RECT 80.295 285.090 80.475 285.445 ;
		LAYER VIA3 ;
		RECT 80.295 288.405 80.475 288.425 ;
		LAYER M1 ;
		RECT 80.295 289.710 80.475 290.105 ;
		LAYER M2 ;
		RECT 80.295 285.755 80.475 285.775 ;
		LAYER M1 ;
		RECT 80.295 288.715 80.475 289.440 ;
		LAYER M2 ;
		RECT 80.295 260.895 80.475 261.580 ;
		LAYER M1 ;
		RECT 80.295 261.870 80.475 262.265 ;
		LAYER M1 ;
		RECT 80.295 262.535 80.475 262.595 ;
		LAYER VIA3 ;
		RECT 80.295 267.855 80.475 268.540 ;
		LAYER VIA3 ;
		RECT 80.295 267.525 80.475 267.545 ;
		LAYER VIA3 ;
		RECT 80.295 265.535 80.475 266.220 ;
		LAYER M2 ;
		RECT 80.295 269.515 80.475 269.535 ;
		LAYER M3 ;
		RECT 80.295 269.515 80.475 269.535 ;
		LAYER VIA3 ;
		RECT 80.295 269.515 80.475 269.535 ;
		LAYER M3 ;
		RECT 80.295 269.845 80.475 269.865 ;
		LAYER M2 ;
		RECT 80.295 270.175 80.475 270.860 ;
		LAYER M3 ;
		RECT 80.295 270.175 80.475 270.860 ;
		LAYER VIA3 ;
		RECT 80.295 270.175 80.475 270.860 ;
		LAYER M1 ;
		RECT 80.295 270.155 80.475 270.880 ;
		LAYER VIA3 ;
		RECT 80.295 272.495 80.475 273.180 ;
		LAYER VIA3 ;
		RECT 80.295 268.850 80.475 269.205 ;
		LAYER VIA3 ;
		RECT 80.295 269.845 80.475 269.865 ;
		LAYER M2 ;
		RECT 80.295 218.805 80.475 218.825 ;
		LAYER M2 ;
		RECT 80.295 218.475 80.475 218.495 ;
		LAYER M1 ;
		RECT 80.295 218.455 80.475 218.515 ;
		LAYER M1 ;
		RECT 80.295 216.465 80.475 216.525 ;
		LAYER M1 ;
		RECT 80.295 206.855 80.475 206.915 ;
		LAYER M1 ;
		RECT 80.295 206.190 80.475 206.585 ;
		LAYER M1 ;
		RECT 80.295 207.185 80.475 207.245 ;
		LAYER M2 ;
		RECT 80.295 213.835 80.475 213.855 ;
		LAYER M3 ;
		RECT 80.295 213.835 80.475 213.855 ;
		LAYER M2 ;
		RECT 80.295 214.165 80.475 214.185 ;
		LAYER M3 ;
		RECT 80.295 214.165 80.475 214.185 ;
		LAYER M3 ;
		RECT 80.295 188.645 80.475 188.665 ;
		LAYER M2 ;
		RECT 80.295 188.645 80.475 188.665 ;
		LAYER M1 ;
		RECT 80.295 184.315 80.475 185.040 ;
		LAYER M1 ;
		RECT 80.295 188.295 80.475 188.355 ;
		LAYER M3 ;
		RECT 80.295 184.335 80.475 185.020 ;
		LAYER VIA3 ;
		RECT 80.295 188.645 80.475 188.665 ;
		LAYER M3 ;
		RECT 80.295 188.315 80.475 188.335 ;
		LAYER M3 ;
		RECT 80.295 187.650 80.475 188.005 ;
		LAYER M2 ;
		RECT 80.295 187.650 80.475 188.005 ;
		LAYER M1 ;
		RECT 80.295 187.630 80.475 188.025 ;
		LAYER M3 ;
		RECT 80.295 181.685 80.475 181.705 ;
		LAYER M1 ;
		RECT 80.295 182.990 80.475 183.385 ;
		LAYER M1 ;
		RECT 80.295 183.655 80.475 183.715 ;
		LAYER M2 ;
		RECT 80.295 184.005 80.475 184.025 ;
		LAYER M2 ;
		RECT 80.295 178.700 80.475 178.725 ;
		LAYER M1 ;
		RECT 80.295 183.985 80.475 184.045 ;
		LAYER M3 ;
		RECT 80.295 188.975 80.475 189.660 ;
		LAYER M1 ;
		RECT 80.295 188.625 80.475 188.685 ;
		LAYER VIA3 ;
		RECT 80.295 188.975 80.475 189.660 ;
		LAYER M2 ;
		RECT 80.295 188.315 80.475 188.335 ;
		LAYER M2 ;
		RECT 80.295 185.330 80.475 185.685 ;
		LAYER M3 ;
		RECT 80.295 186.325 80.475 186.345 ;
		LAYER M3 ;
		RECT 80.295 185.995 80.475 186.015 ;
		LAYER M3 ;
		RECT 80.295 185.330 80.475 185.685 ;
		LAYER M1 ;
		RECT 80.295 190.945 80.475 191.005 ;
		LAYER M3 ;
		RECT 80.295 190.965 80.475 190.985 ;
		LAYER M3 ;
		RECT 80.295 190.635 80.475 190.655 ;
		LAYER M3 ;
		RECT 80.295 189.970 80.475 190.325 ;
		LAYER VIA3 ;
		RECT 80.295 190.965 80.475 190.985 ;
		LAYER M1 ;
		RECT 80.295 195.915 80.475 196.640 ;
		LAYER M3 ;
		RECT 80.295 193.285 80.475 193.305 ;
		LAYER M3 ;
		RECT 80.295 192.955 80.475 192.975 ;
		LAYER M3 ;
		RECT 80.295 192.290 80.475 192.645 ;
		LAYER M3 ;
		RECT 80.295 195.935 80.475 196.620 ;
		LAYER M2 ;
		RECT 80.295 177.710 80.475 178.390 ;
		LAYER M1 ;
		RECT 80.295 188.955 80.475 189.680 ;
		LAYER VIA3 ;
		RECT 80.295 191.295 80.475 191.980 ;
		LAYER M1 ;
		RECT 80.295 191.275 80.475 192.000 ;
		LAYER M1 ;
		RECT 80.295 192.935 80.475 192.995 ;
		LAYER M1 ;
		RECT 80.295 193.265 80.475 193.325 ;
		LAYER M1 ;
		RECT 80.295 193.595 80.475 194.320 ;
		LAYER M1 ;
		RECT 80.295 177.690 80.475 178.410 ;
		LAYER VIA3 ;
		RECT 80.295 177.050 80.475 177.400 ;
		LAYER VIA3 ;
		RECT 80.295 176.720 80.475 176.740 ;
		LAYER M2 ;
		RECT 80.295 175.400 80.475 176.080 ;
		LAYER VIA3 ;
		RECT 80.295 175.070 80.475 175.090 ;
		LAYER VIA3 ;
		RECT 80.295 174.740 80.475 174.760 ;
		LAYER M2 ;
		RECT 80.295 174.410 80.475 174.430 ;
		LAYER M2 ;
		RECT 80.295 173.420 80.475 173.770 ;
		LAYER M3 ;
		RECT 80.295 173.420 80.475 173.770 ;
		LAYER M2 ;
		RECT 80.295 172.430 80.475 173.110 ;
		LAYER M3 ;
		RECT 80.295 172.430 80.475 173.110 ;
		LAYER VIA3 ;
		RECT 80.295 166.850 80.475 166.870 ;
		LAYER M1 ;
		RECT 80.295 162.905 80.475 162.965 ;
		LAYER M2 ;
		RECT 80.295 162.925 80.475 162.945 ;
		LAYER M2 ;
		RECT 80.295 160.045 80.475 161.625 ;
		LAYER M2 ;
		RECT 80.295 159.715 80.475 159.735 ;
		LAYER M1 ;
		RECT 80.295 159.695 80.475 159.755 ;
		LAYER M2 ;
		RECT 80.295 162.265 80.475 162.285 ;
		LAYER M1 ;
		RECT 80.295 156.580 80.475 156.640 ;
		LAYER M1 ;
		RECT 80.295 156.155 80.475 156.310 ;
		LAYER VIA3 ;
		RECT 80.295 143.915 80.475 144.850 ;
		LAYER VIA3 ;
		RECT 80.295 142.265 80.475 142.945 ;
		LAYER VIA3 ;
		RECT 80.295 141.935 80.475 141.955 ;
		LAYER M1 ;
		RECT 80.295 143.235 80.475 143.295 ;
		LAYER M1 ;
		RECT 80.295 142.245 80.475 142.965 ;
		LAYER VIA3 ;
		RECT 80.295 162.595 80.475 162.615 ;
		LAYER M2 ;
		RECT 80.295 162.595 80.475 162.615 ;
		LAYER M1 ;
		RECT 80.295 162.575 80.475 162.635 ;
		LAYER M3 ;
		RECT 80.295 162.925 80.475 162.945 ;
		LAYER M1 ;
		RECT 80.295 20.630 80.475 21.025 ;
		LAYER M2 ;
		RECT 80.295 21.315 80.475 21.335 ;
		LAYER M2 ;
		RECT 80.295 21.645 80.475 21.665 ;
		LAYER M2 ;
		RECT 80.295 21.975 80.475 22.660 ;
		LAYER M3 ;
		RECT 80.295 21.645 80.475 21.665 ;
		LAYER M1 ;
		RECT 80.295 54.435 80.475 55.160 ;
		LAYER M2 ;
		RECT 80.295 53.795 80.475 53.815 ;
		LAYER M1 ;
		RECT 80.295 53.775 80.475 53.835 ;
		LAYER M3 ;
		RECT 80.295 57.770 80.475 58.125 ;
		LAYER M1 ;
		RECT 80.295 55.430 80.475 55.825 ;
		LAYER M2 ;
		RECT 80.295 56.115 80.475 56.135 ;
		LAYER M1 ;
		RECT 80.295 56.425 80.475 56.485 ;
		LAYER M2 ;
		RECT 80.295 55.450 80.475 55.805 ;
		LAYER M2 ;
		RECT 80.295 54.455 80.475 55.140 ;
		LAYER M3 ;
		RECT 80.295 54.455 80.475 55.140 ;
		LAYER VIA3 ;
		RECT 80.295 54.455 80.475 55.140 ;
		LAYER VIA3 ;
		RECT 80.295 54.125 80.475 54.145 ;
		LAYER M2 ;
		RECT 80.295 54.125 80.475 54.145 ;
		LAYER M3 ;
		RECT 80.295 54.125 80.475 54.145 ;
		LAYER VIA3 ;
		RECT 80.295 53.795 80.475 53.815 ;
		LAYER M3 ;
		RECT 80.295 53.795 80.475 53.815 ;
		LAYER M3 ;
		RECT 80.295 63.075 80.475 63.095 ;
		LAYER M1 ;
		RECT 80.295 62.390 80.475 62.785 ;
		LAYER M3 ;
		RECT 80.295 63.735 80.475 64.420 ;
		LAYER VIA3 ;
		RECT 80.295 63.735 80.475 64.420 ;
		LAYER M1 ;
		RECT 80.295 63.385 80.475 63.445 ;
		LAYER M3 ;
		RECT 80.295 60.090 80.475 60.445 ;
		LAYER M1 ;
		RECT 80.295 63.715 80.475 64.440 ;
		LAYER M1 ;
		RECT 80.295 64.710 80.475 65.105 ;
		LAYER VIA3 ;
		RECT 80.295 66.055 80.475 66.740 ;
		LAYER VIA3 ;
		RECT 80.295 65.725 80.475 65.745 ;
		LAYER M1 ;
		RECT 80.295 65.705 80.475 65.765 ;
		LAYER VIA3 ;
		RECT 80.295 60.090 80.475 60.445 ;
		LAYER M3 ;
		RECT 80.295 74.675 80.475 74.695 ;
		LAYER M1 ;
		RECT 80.295 70.345 80.475 70.405 ;
		LAYER VIA3 ;
		RECT 80.295 71.690 80.475 72.045 ;
		LAYER VIA3 ;
		RECT 80.295 72.355 80.475 72.375 ;
		LAYER M2 ;
		RECT 80.295 72.355 80.475 72.375 ;
		LAYER M3 ;
		RECT 80.295 74.010 80.475 74.365 ;
		LAYER M2 ;
		RECT 80.295 67.050 80.475 67.405 ;
		LAYER VIA3 ;
		RECT 80.295 69.370 80.475 69.725 ;
		LAYER M1 ;
		RECT 80.295 70.015 80.475 70.075 ;
		LAYER VIA3 ;
		RECT 80.295 70.365 80.475 70.385 ;
		LAYER M2 ;
		RECT 80.295 62.410 80.475 62.765 ;
		LAYER M3 ;
		RECT 80.295 61.415 80.475 62.100 ;
		LAYER M2 ;
		RECT 80.295 61.415 80.475 62.100 ;
		LAYER M2 ;
		RECT 80.295 61.085 80.475 61.105 ;
		LAYER VIA3 ;
		RECT 80.295 62.410 80.475 62.765 ;
		LAYER M1 ;
		RECT 80.295 61.395 80.475 62.120 ;
		LAYER M2 ;
		RECT 80.295 60.755 80.475 60.775 ;
		LAYER M3 ;
		RECT 80.295 60.755 80.475 60.775 ;
		LAYER VIA3 ;
		RECT 80.295 60.755 80.475 60.775 ;
		LAYER M1 ;
		RECT 80.295 60.735 80.475 60.795 ;
		LAYER M3 ;
		RECT 80.295 61.085 80.475 61.105 ;
		LAYER M2 ;
		RECT 80.295 60.090 80.475 60.445 ;
		LAYER M2 ;
		RECT 80.295 59.095 80.475 59.780 ;
		LAYER M2 ;
		RECT 80.295 58.765 80.475 58.785 ;
		LAYER M3 ;
		RECT 80.295 59.095 80.475 59.780 ;
		LAYER VIA3 ;
		RECT 80.295 59.095 80.475 59.780 ;
		LAYER M1 ;
		RECT 80.295 57.750 80.475 58.145 ;
		LAYER M2 ;
		RECT 80.295 57.770 80.475 58.125 ;
		LAYER M2 ;
		RECT 80.295 58.435 80.475 58.455 ;
		LAYER M3 ;
		RECT 80.295 58.435 80.475 58.455 ;
		LAYER VIA3 ;
		RECT 80.295 58.435 80.475 58.455 ;
		LAYER VIA3 ;
		RECT 80.295 61.085 80.475 61.105 ;
		LAYER M3 ;
		RECT 80.295 58.765 80.475 58.785 ;
		LAYER M1 ;
		RECT 80.295 58.745 80.475 58.805 ;
		LAYER M2 ;
		RECT 80.295 56.775 80.475 57.460 ;
		LAYER M1 ;
		RECT 80.295 56.755 80.475 57.480 ;
		LAYER M2 ;
		RECT 80.295 56.445 80.475 56.465 ;
		LAYER M3 ;
		RECT 80.295 16.675 80.475 16.695 ;
		LAYER M1 ;
		RECT 80.295 19.635 80.475 20.360 ;
		LAYER M1 ;
		RECT 80.295 19.305 80.475 19.365 ;
		LAYER M2 ;
		RECT 80.295 16.675 80.475 16.695 ;
		LAYER VIA3 ;
		RECT 80.295 16.675 80.475 16.695 ;
		LAYER VIA3 ;
		RECT 80.295 18.995 80.475 19.015 ;
		LAYER M2 ;
		RECT 80.295 18.330 80.475 18.685 ;
		LAYER M3 ;
		RECT 80.295 18.330 80.475 18.685 ;
		LAYER VIA3 ;
		RECT 80.295 18.330 80.475 18.685 ;
		LAYER M1 ;
		RECT 80.295 17.315 80.475 18.040 ;
		LAYER M1 ;
		RECT 80.295 18.975 80.475 19.035 ;
		LAYER VIA3 ;
		RECT 80.295 19.325 80.475 19.345 ;
		LAYER M3 ;
		RECT 80.295 19.325 80.475 19.345 ;
		LAYER M3 ;
		RECT 80.295 18.995 80.475 19.015 ;
		LAYER M2 ;
		RECT 80.295 17.335 80.475 18.020 ;
		LAYER M3 ;
		RECT 80.295 17.335 80.475 18.020 ;
		LAYER VIA3 ;
		RECT 80.295 17.335 80.475 18.020 ;
		LAYER M1 ;
		RECT 80.295 16.985 80.475 17.045 ;
		LAYER VIA3 ;
		RECT 80.295 17.005 80.475 17.025 ;
		LAYER M2 ;
		RECT 80.295 19.325 80.475 19.345 ;
		LAYER M2 ;
		RECT 80.295 51.805 80.475 51.825 ;
		LAYER M1 ;
		RECT 80.295 51.785 80.475 51.845 ;
		LAYER VIA3 ;
		RECT 80.295 52.135 80.475 52.820 ;
		LAYER M2 ;
		RECT 80.295 52.135 80.475 52.820 ;
		LAYER M3 ;
		RECT 80.295 51.805 80.475 51.825 ;
		LAYER VIA3 ;
		RECT 80.295 51.805 80.475 51.825 ;
		LAYER M3 ;
		RECT 80.295 52.135 80.475 52.820 ;
		LAYER M1 ;
		RECT 80.295 41.510 80.475 41.905 ;
		LAYER M2 ;
		RECT 80.295 40.535 80.475 41.220 ;
		LAYER VIA3 ;
		RECT 80.295 40.535 80.475 41.220 ;
		LAYER M1 ;
		RECT 80.295 40.515 80.475 41.240 ;
		LAYER M1 ;
		RECT 80.295 39.855 80.475 39.915 ;
		LAYER M2 ;
		RECT 80.295 39.875 80.475 39.895 ;
		LAYER VIA3 ;
		RECT 80.295 39.875 80.475 39.895 ;
		LAYER M2 ;
		RECT 80.295 40.205 80.475 40.225 ;
		LAYER M2 ;
		RECT 80.295 53.130 80.475 53.485 ;
		LAYER M3 ;
		RECT 80.295 53.130 80.475 53.485 ;
		LAYER VIA3 ;
		RECT 80.295 53.130 80.475 53.485 ;
		LAYER M3 ;
		RECT 80.295 51.475 80.475 51.495 ;
		LAYER VIA3 ;
		RECT 80.295 39.210 80.475 39.565 ;
		LAYER VIA3 ;
		RECT 80.295 38.215 80.475 38.900 ;
		LAYER M1 ;
		RECT 80.295 30.905 80.475 30.965 ;
		LAYER M3 ;
		RECT 80.295 30.925 80.475 30.945 ;
		LAYER M3 ;
		RECT 80.295 28.275 80.475 28.295 ;
		LAYER VIA3 ;
		RECT 80.295 28.275 80.475 28.295 ;
		LAYER M2 ;
		RECT 80.295 22.970 80.475 23.325 ;
		LAYER VIA3 ;
		RECT 80.295 22.970 80.475 23.325 ;
		LAYER M1 ;
		RECT 80.295 22.950 80.475 23.345 ;
		LAYER M3 ;
		RECT 80.295 21.975 80.475 22.660 ;
		LAYER VIA3 ;
		RECT 80.295 21.975 80.475 22.660 ;
		LAYER VIA3 ;
		RECT 80.295 21.315 80.475 21.335 ;
		LAYER M1 ;
		RECT 80.295 21.295 80.475 21.355 ;
		LAYER M1 ;
		RECT 80.295 21.955 80.475 22.680 ;
		LAYER VIA3 ;
		RECT 80.295 21.645 80.475 21.665 ;
		LAYER M1 ;
		RECT 80.295 21.625 80.475 21.685 ;
		LAYER M3 ;
		RECT 80.295 21.315 80.475 21.335 ;
		LAYER M2 ;
		RECT 80.295 20.650 80.475 21.005 ;
		LAYER M3 ;
		RECT 80.295 20.650 80.475 21.005 ;
		LAYER M2 ;
		RECT 80.295 19.655 80.475 20.340 ;
		LAYER VIA3 ;
		RECT 80.295 20.650 80.475 21.005 ;
		LAYER VIA3 ;
		RECT 80.295 19.655 80.475 20.340 ;
		LAYER M3 ;
		RECT 80.295 19.655 80.475 20.340 ;
		LAYER M1 ;
		RECT 80.295 48.470 80.475 48.865 ;
		LAYER M3 ;
		RECT 80.295 48.490 80.475 48.845 ;
		LAYER VIA3 ;
		RECT 80.295 48.490 80.475 48.845 ;
		LAYER VIA3 ;
		RECT 80.295 46.835 80.475 46.855 ;
		LAYER M2 ;
		RECT 80.295 46.170 80.475 46.525 ;
		LAYER M3 ;
		RECT 80.295 46.170 80.475 46.525 ;
		LAYER M2 ;
		RECT 80.295 45.175 80.475 45.860 ;
		LAYER M3 ;
		RECT 80.295 45.175 80.475 45.860 ;
		LAYER M1 ;
		RECT 80.295 44.825 80.475 44.885 ;
		LAYER M3 ;
		RECT 80.295 44.845 80.475 44.865 ;
		LAYER VIA3 ;
		RECT 80.295 44.845 80.475 44.865 ;
		LAYER M2 ;
		RECT 80.295 44.515 80.475 44.535 ;
		LAYER M3 ;
		RECT 80.295 44.515 80.475 44.535 ;
		LAYER M3 ;
		RECT 80.295 46.835 80.475 46.855 ;
		LAYER M2 ;
		RECT 80.295 51.475 80.475 51.495 ;
		LAYER M1 ;
		RECT 80.295 51.455 80.475 51.515 ;
		LAYER VIA3 ;
		RECT 80.295 49.155 80.475 49.175 ;
		LAYER M3 ;
		RECT 80.295 49.155 80.475 49.175 ;
		LAYER VIA3 ;
		RECT 80.295 41.530 80.475 41.885 ;
		LAYER VIA3 ;
		RECT 80.295 42.525 80.475 42.545 ;
		LAYER M1 ;
		RECT 80.295 40.185 80.475 40.245 ;
		LAYER M2 ;
		RECT 80.295 41.530 80.475 41.885 ;
		LAYER M1 ;
		RECT 80.295 43.830 80.475 44.225 ;
		LAYER M1 ;
		RECT 80.295 42.505 80.475 42.565 ;
		LAYER M2 ;
		RECT 80.295 42.195 80.475 42.215 ;
		LAYER VIA3 ;
		RECT 80.295 42.195 80.475 42.215 ;
		LAYER M3 ;
		RECT 80.295 42.195 80.475 42.215 ;
		LAYER M2 ;
		RECT 80.295 42.525 80.475 42.545 ;
		LAYER M1 ;
		RECT 80.295 33.555 80.475 34.280 ;
		LAYER VIA3 ;
		RECT 80.295 33.575 80.475 34.260 ;
		LAYER M1 ;
		RECT 80.295 33.225 80.475 33.285 ;
		LAYER M2 ;
		RECT 80.295 33.245 80.475 33.265 ;
		LAYER M3 ;
		RECT 80.295 31.255 80.475 31.940 ;
		LAYER M2 ;
		RECT 80.295 30.925 80.475 30.945 ;
		LAYER VIA3 ;
		RECT 80.295 30.925 80.475 30.945 ;
		LAYER VIA3 ;
		RECT 80.295 32.250 80.475 32.605 ;
		LAYER M2 ;
		RECT 80.295 33.575 80.475 34.260 ;
		LAYER M1 ;
		RECT 80.295 29.910 80.475 30.305 ;
		LAYER M1 ;
		RECT 80.295 28.915 80.475 29.640 ;
		LAYER VIA3 ;
		RECT 80.295 30.595 80.475 30.615 ;
		LAYER M1 ;
		RECT 80.295 30.575 80.475 30.635 ;
		LAYER M2 ;
		RECT 80.295 28.275 80.475 28.295 ;
		LAYER M2 ;
		RECT 80.295 28.605 80.475 28.625 ;
		LAYER M1 ;
		RECT 80.295 28.585 80.475 28.645 ;
		LAYER M2 ;
		RECT 80.295 28.935 80.475 29.620 ;
		LAYER M1 ;
		RECT 80.295 28.255 80.475 28.315 ;
		LAYER VIA3 ;
		RECT 80.295 37.885 80.475 37.905 ;
		LAYER M2 ;
		RECT 80.295 36.890 80.475 37.245 ;
		LAYER M1 ;
		RECT 80.295 35.215 80.475 35.275 ;
		LAYER VIA3 ;
		RECT 80.295 34.570 80.475 34.925 ;
		LAYER M3 ;
		RECT 80.295 34.570 80.475 34.925 ;
		LAYER VIA3 ;
		RECT 80.295 37.555 80.475 37.575 ;
		LAYER M3 ;
		RECT 80.295 37.555 80.475 37.575 ;
		LAYER M2 ;
		RECT 80.295 37.555 80.475 37.575 ;
		LAYER VIA3 ;
		RECT 80.295 36.890 80.475 37.245 ;
		LAYER M3 ;
		RECT 80.295 36.890 80.475 37.245 ;
		LAYER M1 ;
		RECT 80.295 35.875 80.475 36.600 ;
		LAYER M2 ;
		RECT 80.295 35.895 80.475 36.580 ;
		LAYER VIA3 ;
		RECT 80.295 35.895 80.475 36.580 ;
		LAYER M2 ;
		RECT 80.295 35.565 80.475 35.585 ;
		LAYER M1 ;
		RECT 80.295 35.545 80.475 35.605 ;
		LAYER M2 ;
		RECT 80.295 35.235 80.475 35.255 ;
		LAYER M3 ;
		RECT 80.295 35.235 80.475 35.255 ;
		LAYER M3 ;
		RECT 80.295 23.965 80.475 23.985 ;
		LAYER M2 ;
		RECT 80.295 23.965 80.475 23.985 ;
		LAYER VIA3 ;
		RECT 80.295 23.965 80.475 23.985 ;
		LAYER VIA3 ;
		RECT 80.295 23.635 80.475 23.655 ;
		LAYER M2 ;
		RECT 80.295 25.955 80.475 25.975 ;
		LAYER M3 ;
		RECT 80.295 25.955 80.475 25.975 ;
		LAYER VIA3 ;
		RECT 80.295 25.955 80.475 25.975 ;
		LAYER M1 ;
		RECT 80.295 26.595 80.475 27.320 ;
		LAYER M1 ;
		RECT 80.295 26.265 80.475 26.325 ;
		LAYER VIA3 ;
		RECT 80.295 26.285 80.475 26.305 ;
		LAYER M3 ;
		RECT 80.295 24.295 80.475 24.980 ;
		LAYER M2 ;
		RECT 80.295 24.295 80.475 24.980 ;
		LAYER M1 ;
		RECT 80.295 27.590 80.475 27.985 ;
		LAYER VIA3 ;
		RECT 80.295 24.295 80.475 24.980 ;
		LAYER M3 ;
		RECT 80.295 25.290 80.475 25.645 ;
		LAYER M2 ;
		RECT 80.295 25.290 80.475 25.645 ;
		LAYER VIA3 ;
		RECT 80.295 25.290 80.475 25.645 ;
		LAYER M1 ;
		RECT 80.295 25.935 80.475 25.995 ;
		LAYER M1 ;
		RECT 80.295 47.475 80.475 48.200 ;
		LAYER M2 ;
		RECT 80.295 47.165 80.475 47.185 ;
		LAYER M3 ;
		RECT 80.295 47.165 80.475 47.185 ;
		LAYER VIA3 ;
		RECT 80.295 47.165 80.475 47.185 ;
		LAYER M2 ;
		RECT 80.295 47.495 80.475 48.180 ;
		LAYER M3 ;
		RECT 80.295 47.495 80.475 48.180 ;
		LAYER VIA3 ;
		RECT 80.295 47.495 80.475 48.180 ;
		LAYER M1 ;
		RECT 80.295 42.835 80.475 43.560 ;
		LAYER M2 ;
		RECT 80.295 43.850 80.475 44.205 ;
		LAYER M3 ;
		RECT 80.295 43.850 80.475 44.205 ;
		LAYER VIA3 ;
		RECT 80.295 43.850 80.475 44.205 ;
		LAYER VIA3 ;
		RECT 80.295 45.175 80.475 45.860 ;
		LAYER M1 ;
		RECT 80.295 216.135 80.475 216.195 ;
		LAYER M2 ;
		RECT 80.295 216.155 80.475 216.175 ;
		LAYER M3 ;
		RECT 80.295 216.155 80.475 216.175 ;
		LAYER M2 ;
		RECT 80.295 213.170 80.475 213.525 ;
		LAYER M1 ;
		RECT 80.295 215.470 80.475 215.865 ;
		LAYER M2 ;
		RECT 80.295 214.495 80.475 215.180 ;
		LAYER M3 ;
		RECT 80.295 214.495 80.475 215.180 ;
		LAYER M2 ;
		RECT 80.295 215.490 80.475 215.845 ;
		LAYER M3 ;
		RECT 80.295 215.490 80.475 215.845 ;
		LAYER VIA3 ;
		RECT 80.295 214.495 80.475 215.180 ;
		LAYER M2 ;
		RECT 80.295 212.175 80.475 212.860 ;
		LAYER M3 ;
		RECT 80.295 212.175 80.475 212.860 ;
		LAYER M2 ;
		RECT 80.295 211.845 80.475 211.865 ;
		LAYER M3 ;
		RECT 80.295 211.845 80.475 211.865 ;
		LAYER M2 ;
		RECT 80.295 210.850 80.475 211.205 ;
		LAYER M3 ;
		RECT 80.295 210.850 80.475 211.205 ;
		LAYER M2 ;
		RECT 80.295 211.515 80.475 211.535 ;
		LAYER M3 ;
		RECT 80.295 211.515 80.475 211.535 ;
		LAYER VIA3 ;
		RECT 80.295 211.515 80.475 211.535 ;
		LAYER M1 ;
		RECT 80.295 209.505 80.475 209.565 ;
		LAYER M1 ;
		RECT 80.295 209.175 80.475 209.235 ;
		LAYER M3 ;
		RECT 80.295 213.170 80.475 213.525 ;
		LAYER M3 ;
		RECT 80.295 209.855 80.475 210.540 ;
		LAYER VIA3 ;
		RECT 80.295 209.855 80.475 210.540 ;
		LAYER M2 ;
		RECT 80.295 171.110 80.475 171.130 ;
		LAYER M3 ;
		RECT 80.295 171.110 80.475 171.130 ;
		LAYER VIA3 ;
		RECT 80.295 171.440 80.475 171.460 ;
		LAYER M1 ;
		RECT 80.295 171.420 80.475 171.480 ;
		LAYER M2 ;
		RECT 80.295 171.440 80.475 171.460 ;
		LAYER VIA3 ;
		RECT 80.295 171.110 80.475 171.130 ;
		LAYER VIA3 ;
		RECT 80.295 174.410 80.475 174.430 ;
		LAYER M1 ;
		RECT 80.295 174.390 80.475 174.450 ;
		LAYER M2 ;
		RECT 80.295 174.740 80.475 174.760 ;
		LAYER M2 ;
		RECT 80.295 175.070 80.475 175.090 ;
		LAYER M1 ;
		RECT 80.295 174.720 80.475 174.780 ;
		LAYER M2 ;
		RECT 80.295 171.770 80.475 172.120 ;
		LAYER M2 ;
		RECT 80.295 176.390 80.475 176.410 ;
		LAYER M1 ;
		RECT 80.295 175.050 80.475 175.110 ;
		LAYER M1 ;
		RECT 80.295 171.750 80.475 172.140 ;
		LAYER M1 ;
		RECT 80.295 177.030 80.475 177.420 ;
		LAYER M1 ;
		RECT 80.295 176.700 80.475 176.760 ;
		LAYER M3 ;
		RECT 80.295 177.710 80.475 178.390 ;
		LAYER M3 ;
		RECT 80.295 178.700 80.475 178.725 ;
		LAYER M1 ;
		RECT 80.295 205.195 80.475 205.920 ;
		LAYER M2 ;
		RECT 80.295 204.885 80.475 204.905 ;
		LAYER M3 ;
		RECT 80.295 204.885 80.475 204.905 ;
		LAYER VIA3 ;
		RECT 80.295 204.885 80.475 204.905 ;
		LAYER M2 ;
		RECT 80.295 170.120 80.475 170.800 ;
		LAYER VIA3 ;
		RECT 80.295 170.120 80.475 170.800 ;
		LAYER M1 ;
		RECT 80.295 198.235 80.475 198.960 ;
		LAYER M1 ;
		RECT 80.295 171.090 80.475 171.150 ;
		LAYER VIA3 ;
		RECT 80.295 197.925 80.475 197.945 ;
		LAYER M1 ;
		RECT 80.295 197.905 80.475 197.965 ;
		LAYER M1 ;
		RECT 80.295 202.875 80.475 203.600 ;
		LAYER VIA3 ;
		RECT 80.295 202.895 80.475 203.580 ;
		LAYER VIA3 ;
		RECT 80.295 202.235 80.475 202.255 ;
		LAYER M2 ;
		RECT 80.295 199.250 80.475 199.605 ;
		LAYER M1 ;
		RECT 80.295 200.225 80.475 200.285 ;
		LAYER VIA3 ;
		RECT 80.295 200.245 80.475 200.265 ;
		LAYER M2 ;
		RECT 80.295 200.245 80.475 200.265 ;
		LAYER M1 ;
		RECT 80.295 199.895 80.475 199.955 ;
		LAYER M3 ;
		RECT 80.295 200.245 80.475 200.265 ;
		LAYER M1 ;
		RECT 80.295 199.230 80.475 199.625 ;
		LAYER M2 ;
		RECT 80.295 199.915 80.475 199.935 ;
		LAYER M3 ;
		RECT 80.295 199.915 80.475 199.935 ;
		LAYER VIA3 ;
		RECT 80.295 199.915 80.475 199.935 ;
		LAYER VIA3 ;
		RECT 80.295 199.250 80.475 199.605 ;
		LAYER M3 ;
		RECT 80.295 199.250 80.475 199.605 ;
		LAYER M2 ;
		RECT 80.295 200.575 80.475 201.260 ;
		LAYER M1 ;
		RECT 80.295 200.555 80.475 201.280 ;
		LAYER VIA3 ;
		RECT 80.295 201.570 80.475 201.925 ;
		LAYER M3 ;
		RECT 80.295 198.255 80.475 198.940 ;
		LAYER M2 ;
		RECT 80.295 202.565 80.475 202.585 ;
		LAYER VIA3 ;
		RECT 80.295 202.565 80.475 202.585 ;
		LAYER M1 ;
		RECT 80.295 202.545 80.475 202.605 ;
		LAYER M2 ;
		RECT 80.295 202.235 80.475 202.255 ;
		LAYER M3 ;
		RECT 80.295 202.235 80.475 202.255 ;
		LAYER M3 ;
		RECT 80.295 202.565 80.475 202.585 ;
		LAYER VIA3 ;
		RECT 80.295 200.575 80.475 201.260 ;
		LAYER VIA3 ;
		RECT 80.295 198.255 80.475 198.940 ;
		LAYER M2 ;
		RECT 80.295 198.255 80.475 198.940 ;
		LAYER M3 ;
		RECT 80.295 200.575 80.475 201.260 ;
		LAYER M3 ;
		RECT 80.295 171.770 80.475 172.120 ;
		LAYER M2 ;
		RECT 80.295 176.720 80.475 176.740 ;
		LAYER M3 ;
		RECT 80.295 176.720 80.475 176.740 ;
		LAYER M1 ;
		RECT 80.295 179.015 80.475 179.075 ;
		LAYER M3 ;
		RECT 80.295 177.050 80.475 177.400 ;
		LAYER M3 ;
		RECT 80.295 174.410 80.475 174.430 ;
		LAYER M3 ;
		RECT 80.295 174.080 80.475 174.100 ;
		LAYER M3 ;
		RECT 80.295 175.400 80.475 176.080 ;
		LAYER VIA3 ;
		RECT 80.295 175.400 80.475 176.080 ;
		LAYER M3 ;
		RECT 80.295 183.675 80.475 183.695 ;
		LAYER M3 ;
		RECT 80.295 184.005 80.475 184.025 ;
		LAYER M2 ;
		RECT 80.295 184.335 80.475 185.020 ;
		LAYER M2 ;
		RECT 80.295 185.995 80.475 186.015 ;
		LAYER M1 ;
		RECT 80.295 175.380 80.475 176.100 ;
		LAYER M3 ;
		RECT 80.295 176.390 80.475 176.410 ;
		LAYER VIA3 ;
		RECT 80.295 176.390 80.475 176.410 ;
		LAYER M1 ;
		RECT 80.295 176.370 80.475 176.430 ;
		LAYER M2 ;
		RECT 80.295 179.035 80.475 179.055 ;
		LAYER M2 ;
		RECT 80.295 179.365 80.475 179.385 ;
		LAYER VIA3 ;
		RECT 80.295 179.365 80.475 179.385 ;
		LAYER M3 ;
		RECT 80.295 179.365 80.475 179.385 ;
		LAYER VIA3 ;
		RECT 80.295 179.035 80.475 179.055 ;
		LAYER M3 ;
		RECT 80.295 179.035 80.475 179.055 ;
		LAYER M1 ;
		RECT 80.295 179.345 80.475 179.405 ;
		LAYER M1 ;
		RECT 80.295 181.995 80.475 182.720 ;
		LAYER VIA3 ;
		RECT 80.295 185.995 80.475 186.015 ;
		LAYER M1 ;
		RECT 80.295 185.310 80.475 185.705 ;
		LAYER M1 ;
		RECT 80.295 218.785 80.475 218.845 ;
		LAYER VIA3 ;
		RECT 80.295 117.095 80.475 117.780 ;
		LAYER M3 ;
		RECT 80.295 160.045 80.475 161.625 ;
		LAYER VIA3 ;
		RECT 80.295 157.815 80.475 159.405 ;
		LAYER M3 ;
		RECT 80.295 157.815 80.475 159.405 ;
		LAYER M2 ;
		RECT 80.295 157.815 80.475 159.405 ;
		LAYER M2 ;
		RECT 80.295 216.815 80.475 217.500 ;
		LAYER M2 ;
		RECT 80.295 161.935 80.475 161.955 ;
		LAYER VIA3 ;
		RECT 80.295 161.935 80.475 161.955 ;
		LAYER M1 ;
		RECT 80.295 164.850 80.475 166.230 ;
		LAYER M2 ;
		RECT 80.295 217.810 80.475 218.165 ;
		LAYER VIA3 ;
		RECT 80.295 160.045 80.475 161.625 ;
		LAYER M3 ;
		RECT 80.295 161.935 80.475 161.955 ;
		LAYER M1 ;
		RECT 80.295 161.915 80.475 161.975 ;
		LAYER M2 ;
		RECT 80.295 166.850 80.475 166.870 ;
		LAYER VIA3 ;
		RECT 80.295 164.870 80.475 166.210 ;
		LAYER M3 ;
		RECT 80.295 164.870 80.475 166.210 ;
		LAYER M2 ;
		RECT 80.295 157.485 80.475 157.505 ;
		LAYER M3 ;
		RECT 80.295 156.930 80.475 157.175 ;
		LAYER M1 ;
		RECT 80.295 156.910 80.475 157.195 ;
		LAYER VIA3 ;
		RECT 80.295 157.485 80.475 157.505 ;
		LAYER M3 ;
		RECT 80.295 157.485 80.475 157.505 ;
		LAYER VIA3 ;
		RECT 80.295 156.930 80.475 157.175 ;
		LAYER VIA3 ;
		RECT 80.295 156.175 80.475 156.290 ;
		LAYER M2 ;
		RECT 80.295 156.175 80.475 156.290 ;
		LAYER M3 ;
		RECT 80.295 156.175 80.475 156.290 ;
		LAYER VIA3 ;
		RECT 80.295 155.015 80.475 155.865 ;
		LAYER M2 ;
		RECT 80.295 155.015 80.475 155.865 ;
		LAYER M3 ;
		RECT 80.295 155.015 80.475 155.865 ;
		LAYER M1 ;
		RECT 80.295 154.995 80.475 155.885 ;
		LAYER M2 ;
		RECT 80.295 140.285 80.475 140.965 ;
		LAYER M3 ;
		RECT 80.295 140.285 80.475 140.965 ;
		LAYER M1 ;
		RECT 80.295 140.265 80.475 140.985 ;
		LAYER M3 ;
		RECT 80.295 141.275 80.475 141.295 ;
		LAYER M2 ;
		RECT 80.295 138.965 80.475 138.985 ;
		LAYER M3 ;
		RECT 80.295 138.965 80.475 138.985 ;
		LAYER VIA3 ;
		RECT 80.295 138.965 80.475 138.985 ;
		LAYER M1 ;
		RECT 80.295 138.945 80.475 139.005 ;
		LAYER M3 ;
		RECT 80.295 139.295 80.475 139.315 ;
		LAYER M1 ;
		RECT 80.295 137.955 80.475 138.675 ;
		LAYER VIA3 ;
		RECT 80.295 137.975 80.475 138.655 ;
		LAYER M3 ;
		RECT 80.295 146.810 80.475 146.830 ;
		LAYER VIA3 ;
		RECT 80.295 146.810 80.475 146.830 ;
		LAYER M1 ;
		RECT 80.295 146.460 80.475 146.520 ;
		LAYER M3 ;
		RECT 80.295 141.935 80.475 141.955 ;
		LAYER M1 ;
		RECT 80.295 141.255 80.475 141.315 ;
		LAYER M2 ;
		RECT 80.295 141.275 80.475 141.295 ;
		LAYER M1 ;
		RECT 80.295 141.585 80.475 141.645 ;
		LAYER M2 ;
		RECT 80.295 153.285 80.475 153.305 ;
		LAYER VIA3 ;
		RECT 80.295 153.285 80.475 153.305 ;
		LAYER M3 ;
		RECT 80.295 154.305 80.475 154.705 ;
		LAYER M1 ;
		RECT 80.295 153.595 80.475 153.685 ;
		LAYER M1 ;
		RECT 80.295 153.265 80.475 153.325 ;
		LAYER M3 ;
		RECT 80.295 153.285 80.475 153.305 ;
		LAYER VIA3 ;
		RECT 80.295 152.495 80.475 152.975 ;
		LAYER M3 ;
		RECT 80.295 148.855 80.475 148.875 ;
		LAYER M1 ;
		RECT 80.295 152.475 80.475 152.995 ;
		LAYER VIA3 ;
		RECT 80.295 152.165 80.475 152.185 ;
		LAYER M3 ;
		RECT 80.295 152.165 80.475 152.185 ;
		LAYER VIA3 ;
		RECT 80.295 149.185 80.475 151.855 ;
		LAYER VIA3 ;
		RECT 80.295 148.855 80.475 148.875 ;
		LAYER M1 ;
		RECT 80.295 148.835 80.475 148.895 ;
		LAYER VIA3 ;
		RECT 80.295 139.295 80.475 139.315 ;
		LAYER M3 ;
		RECT 80.295 147.140 80.475 147.840 ;
		LAYER M1 ;
		RECT 80.295 148.130 80.475 148.235 ;
		LAYER M1 ;
		RECT 80.295 147.120 80.475 147.860 ;
		LAYER VIA3 ;
		RECT 80.295 153.615 80.475 153.665 ;
		LAYER M2 ;
		RECT 80.295 153.615 80.475 153.665 ;
		LAYER M2 ;
		RECT 80.295 154.305 80.475 154.705 ;
		LAYER M3 ;
		RECT 80.295 153.615 80.475 153.665 ;
		LAYER VIA3 ;
		RECT 80.295 153.975 80.475 153.995 ;
		LAYER M2 ;
		RECT 80.295 153.975 80.475 153.995 ;
		LAYER M1 ;
		RECT 80.295 153.955 80.475 154.015 ;
		LAYER VIA3 ;
		RECT 80.295 154.305 80.475 154.705 ;
		LAYER M2 ;
		RECT 80.295 141.605 80.475 141.625 ;
		LAYER M3 ;
		RECT 80.295 141.605 80.475 141.625 ;
		LAYER VIA3 ;
		RECT 80.295 141.605 80.475 141.625 ;
		LAYER M2 ;
		RECT 80.295 141.935 80.475 141.955 ;
		LAYER M2 ;
		RECT 80.295 142.265 80.475 142.945 ;
		LAYER M3 ;
		RECT 80.295 146.150 80.475 146.170 ;
		LAYER M1 ;
		RECT 80.295 145.140 80.475 145.860 ;
		LAYER M1 ;
		RECT 80.295 143.895 80.475 144.870 ;
		LAYER M2 ;
		RECT 80.295 146.810 80.475 146.830 ;
		LAYER M1 ;
		RECT 80.295 146.790 80.475 146.850 ;
		LAYER VIA3 ;
		RECT 80.295 146.480 80.475 146.500 ;
		LAYER M2 ;
		RECT 80.295 146.480 80.475 146.500 ;
		LAYER M3 ;
		RECT 80.295 146.480 80.475 146.500 ;
		LAYER M2 ;
		RECT 80.295 147.140 80.475 147.840 ;
		LAYER VIA3 ;
		RECT 80.295 147.140 80.475 147.840 ;
		LAYER VIA3 ;
		RECT 80.295 146.150 80.475 146.170 ;
		LAYER M2 ;
		RECT 80.295 146.150 80.475 146.170 ;
		LAYER M2 ;
		RECT 80.295 156.930 80.475 157.175 ;
		LAYER VIA3 ;
		RECT 80.295 133.335 80.475 134.020 ;
		LAYER M1 ;
		RECT 80.295 129.670 80.475 130.065 ;
		LAYER M1 ;
		RECT 80.295 128.675 80.475 129.400 ;
		LAYER M1 ;
		RECT 80.295 154.285 80.475 154.725 ;
		LAYER M1 ;
		RECT 80.295 164.520 80.475 164.580 ;
		LAYER M3 ;
		RECT 80.295 164.540 80.475 164.560 ;
		LAYER M3 ;
		RECT 80.295 164.210 80.475 164.230 ;
		LAYER M2 ;
		RECT 80.295 164.210 80.475 164.230 ;
		LAYER M2 ;
		RECT 80.295 164.540 80.475 164.560 ;
		LAYER M1 ;
		RECT 80.295 163.235 80.475 163.295 ;
		LAYER M3 ;
		RECT 80.295 159.715 80.475 159.735 ;
		LAYER VIA3 ;
		RECT 80.295 159.715 80.475 159.735 ;
		LAYER VIA3 ;
		RECT 80.295 162.925 80.475 162.945 ;
		LAYER VIA3 ;
		RECT 80.295 162.265 80.475 162.285 ;
		LAYER M3 ;
		RECT 80.295 162.265 80.475 162.285 ;
		LAYER M1 ;
		RECT 80.295 162.245 80.475 162.305 ;
		LAYER M3 ;
		RECT 80.295 79.315 80.475 79.335 ;
		LAYER M3 ;
		RECT 80.295 86.935 80.475 87.620 ;
		LAYER M1 ;
		RECT 80.295 90.895 80.475 90.955 ;
		LAYER VIA3 ;
		RECT 80.295 82.295 80.475 82.980 ;
		LAYER M3 ;
		RECT 80.295 82.295 80.475 82.980 ;
		LAYER M1 ;
		RECT 80.295 81.945 80.475 82.005 ;
		LAYER M3 ;
		RECT 80.295 81.635 80.475 81.655 ;
		LAYER VIA3 ;
		RECT 80.295 97.875 80.475 97.895 ;
		LAYER M1 ;
		RECT 80.295 97.855 80.475 97.915 ;
		LAYER M1 ;
		RECT 80.295 97.190 80.475 97.585 ;
		LAYER M2 ;
		RECT 80.295 97.875 80.475 97.895 ;
		LAYER M3 ;
		RECT 80.295 97.875 80.475 97.895 ;
		LAYER VIA3 ;
		RECT 80.295 84.285 80.475 84.305 ;
		LAYER VIA3 ;
		RECT 80.295 83.955 80.475 83.975 ;
		LAYER VIA3 ;
		RECT 80.295 85.610 80.475 85.965 ;
		LAYER M1 ;
		RECT 80.295 86.585 80.475 86.645 ;
		LAYER M1 ;
		RECT 80.295 96.195 80.475 96.920 ;
		LAYER M2 ;
		RECT 80.295 90.915 80.475 90.935 ;
		LAYER M3 ;
		RECT 80.295 90.915 80.475 90.935 ;
		LAYER M1 ;
		RECT 80.295 91.225 80.475 91.285 ;
		LAYER M1 ;
		RECT 80.295 95.865 80.475 95.925 ;
		LAYER M1 ;
		RECT 80.295 95.535 80.475 95.595 ;
		LAYER M3 ;
		RECT 80.295 93.895 80.475 94.580 ;
		LAYER M1 ;
		RECT 80.295 93.545 80.475 93.605 ;
		LAYER M2 ;
		RECT 80.295 92.570 80.475 92.925 ;
		LAYER VIA3 ;
		RECT 80.295 91.575 80.475 92.260 ;
		LAYER M1 ;
		RECT 80.295 91.555 80.475 92.280 ;
		LAYER M3 ;
		RECT 80.295 91.245 80.475 91.265 ;
		LAYER VIA3 ;
		RECT 80.295 97.210 80.475 97.565 ;
		LAYER M2 ;
		RECT 80.295 97.210 80.475 97.565 ;
		LAYER M3 ;
		RECT 80.295 97.210 80.475 97.565 ;
		LAYER VIA3 ;
		RECT 80.295 96.215 80.475 96.900 ;
		LAYER VIA3 ;
		RECT 80.295 106.490 80.475 106.845 ;
		LAYER M2 ;
		RECT 80.295 106.490 80.475 106.845 ;
		LAYER M3 ;
		RECT 80.295 106.490 80.475 106.845 ;
		LAYER M1 ;
		RECT 80.295 106.470 80.475 106.865 ;
		LAYER VIA3 ;
		RECT 80.295 107.155 80.475 107.175 ;
		LAYER M2 ;
		RECT 80.295 107.155 80.475 107.175 ;
		LAYER M3 ;
		RECT 80.295 107.155 80.475 107.175 ;
		LAYER M2 ;
		RECT 80.295 107.815 80.475 108.500 ;
		LAYER M2 ;
		RECT 80.295 107.485 80.475 107.505 ;
		LAYER M3 ;
		RECT 80.295 107.485 80.475 107.505 ;
		LAYER VIA3 ;
		RECT 80.295 107.485 80.475 107.505 ;
		LAYER M3 ;
		RECT 80.295 107.815 80.475 108.500 ;
		LAYER VIA3 ;
		RECT 80.295 107.815 80.475 108.500 ;
		LAYER M1 ;
		RECT 80.295 107.465 80.475 107.525 ;
		LAYER VIA3 ;
		RECT 80.295 68.375 80.475 69.060 ;
		LAYER VIA3 ;
		RECT 80.295 68.045 80.475 68.065 ;
		LAYER M3 ;
		RECT 80.295 67.050 80.475 67.405 ;
		LAYER M1 ;
		RECT 80.295 67.030 80.475 67.425 ;
		LAYER VIA3 ;
		RECT 80.295 67.050 80.475 67.405 ;
		LAYER VIA3 ;
		RECT 80.295 70.695 80.475 71.380 ;
		LAYER M1 ;
		RECT 80.295 53.110 80.475 53.505 ;
		LAYER M1 ;
		RECT 80.295 52.115 80.475 52.840 ;
		LAYER M1 ;
		RECT 80.295 46.150 80.475 46.545 ;
		LAYER M1 ;
		RECT 80.295 45.155 80.475 45.880 ;
		LAYER M3 ;
		RECT 80.295 37.885 80.475 37.905 ;
		LAYER M2 ;
		RECT 80.295 37.885 80.475 37.905 ;
		LAYER M2 ;
		RECT 80.295 38.215 80.475 38.900 ;
		LAYER M2 ;
		RECT 80.295 39.210 80.475 39.565 ;
		LAYER M3 ;
		RECT 80.295 33.245 80.475 33.265 ;
		LAYER VIA3 ;
		RECT 80.295 33.245 80.475 33.265 ;
		LAYER M3 ;
		RECT 80.295 32.915 80.475 32.935 ;
		LAYER M2 ;
		RECT 80.295 32.250 80.475 32.605 ;
		LAYER M3 ;
		RECT 80.295 35.895 80.475 36.580 ;
		LAYER M3 ;
		RECT 80.295 35.565 80.475 35.585 ;
		LAYER M1 ;
		RECT 80.295 36.870 80.475 37.265 ;
		LAYER M1 ;
		RECT 80.295 34.550 80.475 34.945 ;
		LAYER M2 ;
		RECT 80.295 34.570 80.475 34.925 ;
		LAYER M2 ;
		RECT 80.295 63.405 80.475 63.425 ;
		LAYER M3 ;
		RECT 80.295 63.405 80.475 63.425 ;
		LAYER M1 ;
		RECT 80.295 60.070 80.475 60.465 ;
		LAYER M1 ;
		RECT 80.295 59.075 80.475 59.800 ;
		LAYER VIA3 ;
		RECT 80.295 72.685 80.475 72.705 ;
		LAYER M2 ;
		RECT 80.295 72.685 80.475 72.705 ;
		LAYER M3 ;
		RECT 80.295 72.355 80.475 72.375 ;
		LAYER M3 ;
		RECT 80.295 72.685 80.475 72.705 ;
		LAYER M1 ;
		RECT 80.295 73.990 80.475 74.385 ;
		LAYER M2 ;
		RECT 80.295 74.010 80.475 74.365 ;
		LAYER M3 ;
		RECT 80.295 73.015 80.475 73.700 ;
		LAYER M1 ;
		RECT 80.295 72.995 80.475 73.720 ;
		LAYER VIA3 ;
		RECT 80.295 74.675 80.475 74.695 ;
		LAYER M1 ;
		RECT 80.295 74.655 80.475 74.715 ;
		LAYER VIA3 ;
		RECT 80.295 75.005 80.475 75.025 ;
		LAYER M2 ;
		RECT 80.295 75.005 80.475 75.025 ;
		LAYER VIA3 ;
		RECT 80.295 92.570 80.475 92.925 ;
		LAYER M2 ;
		RECT 80.295 84.615 80.475 85.300 ;
		LAYER M2 ;
		RECT 80.295 84.285 80.475 84.305 ;
		LAYER M3 ;
		RECT 80.295 84.285 80.475 84.305 ;
		LAYER M3 ;
		RECT 80.295 83.955 80.475 83.975 ;
		LAYER M1 ;
		RECT 80.295 89.235 80.475 89.960 ;
		LAYER M2 ;
		RECT 80.295 74.675 80.475 74.695 ;
		LAYER M2 ;
		RECT 80.295 79.975 80.475 80.660 ;
		LAYER M3 ;
		RECT 80.295 79.975 80.475 80.660 ;
		LAYER M2 ;
		RECT 80.295 75.335 80.475 76.020 ;
		LAYER M2 ;
		RECT 80.295 77.655 80.475 78.340 ;
		LAYER M3 ;
		RECT 80.295 77.655 80.475 78.340 ;
		LAYER M2 ;
		RECT 80.295 79.645 80.475 79.665 ;
		LAYER M3 ;
		RECT 80.295 79.645 80.475 79.665 ;
		LAYER M3 ;
		RECT 80.295 64.730 80.475 65.085 ;
		LAYER M2 ;
		RECT 80.295 65.395 80.475 65.415 ;
		LAYER M3 ;
		RECT 80.295 65.395 80.475 65.415 ;
		LAYER M1 ;
		RECT 80.295 65.375 80.475 65.435 ;
		LAYER M2 ;
		RECT 80.295 64.730 80.475 65.085 ;
		LAYER M1 ;
		RECT 80.295 92.550 80.475 92.945 ;
		LAYER M2 ;
		RECT 80.295 91.575 80.475 92.260 ;
		LAYER M2 ;
		RECT 80.295 91.245 80.475 91.265 ;
		LAYER M1 ;
		RECT 80.295 90.230 80.475 90.625 ;
		LAYER VIA3 ;
		RECT 80.295 95.885 80.475 95.905 ;
		LAYER VIA3 ;
		RECT 80.295 95.555 80.475 95.575 ;
		LAYER VIA3 ;
		RECT 80.295 94.890 80.475 95.245 ;
		LAYER VIA3 ;
		RECT 80.295 93.235 80.475 93.255 ;
		LAYER VIA3 ;
		RECT 80.295 93.895 80.475 94.580 ;
		LAYER M3 ;
		RECT 80.295 96.215 80.475 96.900 ;
		LAYER M1 ;
		RECT 80.295 113.430 80.475 113.825 ;
		LAYER M2 ;
		RECT 80.295 113.450 80.475 113.805 ;
		LAYER M2 ;
		RECT 80.295 114.115 80.475 114.135 ;
		LAYER M3 ;
		RECT 80.295 114.115 80.475 114.135 ;
		LAYER VIA3 ;
		RECT 80.295 114.115 80.475 114.135 ;
		LAYER VIA3 ;
		RECT 80.295 109.475 80.475 109.495 ;
		LAYER M1 ;
		RECT 80.295 109.455 80.475 109.515 ;
		LAYER M2 ;
		RECT 80.295 109.805 80.475 109.825 ;
		LAYER VIA3 ;
		RECT 80.295 109.805 80.475 109.825 ;
		LAYER VIA3 ;
		RECT 80.295 108.810 80.475 109.165 ;
		LAYER M2 ;
		RECT 80.295 111.130 80.475 111.485 ;
		LAYER M1 ;
		RECT 80.295 111.110 80.475 111.505 ;
		LAYER VIA3 ;
		RECT 80.295 111.130 80.475 111.485 ;
		LAYER M2 ;
		RECT 80.295 265.205 80.475 265.225 ;
		LAYER M1 ;
		RECT 80.295 265.185 80.475 265.245 ;
		LAYER M3 ;
		RECT 80.295 263.215 80.475 263.900 ;
		LAYER M1 ;
		RECT 80.295 264.855 80.475 264.915 ;
		LAYER VIA3 ;
		RECT 80.295 264.210 80.475 264.565 ;
		LAYER M1 ;
		RECT 80.295 264.190 80.475 264.585 ;
		LAYER M2 ;
		RECT 80.295 263.215 80.475 263.900 ;
		LAYER VIA3 ;
		RECT 80.295 263.215 80.475 263.900 ;
		LAYER M1 ;
		RECT 80.295 263.195 80.475 263.920 ;
		LAYER VIA3 ;
		RECT 80.295 239.685 80.475 239.705 ;
		LAYER M3 ;
		RECT 80.295 238.690 80.475 239.045 ;
		LAYER M3 ;
		RECT 80.295 230.405 80.475 230.425 ;
		LAYER M3 ;
		RECT 80.295 230.735 80.475 231.420 ;
		LAYER M3 ;
		RECT 80.295 232.395 80.475 232.415 ;
		LAYER VIA3 ;
		RECT 80.295 232.725 80.475 232.745 ;
		LAYER M2 ;
		RECT 80.295 262.885 80.475 262.905 ;
		LAYER M3 ;
		RECT 80.295 262.885 80.475 262.905 ;
		LAYER VIA3 ;
		RECT 80.295 244.655 80.475 245.340 ;
		LAYER M1 ;
		RECT 80.295 244.305 80.475 244.365 ;
		LAYER M2 ;
		RECT 80.295 244.655 80.475 245.340 ;
		LAYER M3 ;
		RECT 80.295 244.655 80.475 245.340 ;
		LAYER M3 ;
		RECT 80.295 230.075 80.475 230.095 ;
		LAYER M3 ;
		RECT 80.295 228.415 80.475 229.100 ;
		LAYER VIA3 ;
		RECT 80.295 233.055 80.475 233.740 ;
		LAYER M3 ;
		RECT 80.295 3.085 80.475 3.105 ;
		LAYER VIA3 ;
		RECT 80.295 14.685 80.475 14.705 ;
		LAYER M1 ;
		RECT 80.295 14.335 80.475 14.395 ;
		LAYER M1 ;
		RECT 80.295 3.395 80.475 4.120 ;
		LAYER M2 ;
		RECT 80.295 3.085 80.475 3.105 ;
		LAYER VIA3 ;
		RECT 80.295 3.085 80.475 3.105 ;
		LAYER M2 ;
		RECT 80.295 3.415 80.475 4.100 ;
		LAYER M1 ;
		RECT 80.295 12.675 80.475 13.400 ;
		LAYER M1 ;
		RECT 80.295 4.390 80.475 4.785 ;
		LAYER M3 ;
		RECT 80.295 3.415 80.475 4.100 ;
		LAYER VIA3 ;
		RECT 80.295 3.415 80.475 4.100 ;
		LAYER M3 ;
		RECT 80.295 12.365 80.475 12.385 ;
		LAYER VIA3 ;
		RECT 80.295 12.365 80.475 12.385 ;
		LAYER M2 ;
		RECT 80.295 12.365 80.475 12.385 ;
		LAYER M1 ;
		RECT 80.295 12.345 80.475 12.405 ;
		LAYER M3 ;
		RECT 80.295 14.685 80.475 14.705 ;
		LAYER M2 ;
		RECT 80.295 14.685 80.475 14.705 ;
		LAYER VIA3 ;
		RECT 80.295 15.015 80.475 15.700 ;
		LAYER M3 ;
		RECT 80.295 15.015 80.475 15.700 ;
		LAYER M2 ;
		RECT 80.295 4.410 80.475 4.765 ;
		LAYER M1 ;
		RECT 80.295 10.355 80.475 11.080 ;
		LAYER M1 ;
		RECT 80.295 5.055 80.475 5.115 ;
		LAYER M3 ;
		RECT 80.295 4.410 80.475 4.765 ;
		LAYER VIA3 ;
		RECT 80.295 4.410 80.475 4.765 ;
		LAYER M3 ;
		RECT 80.295 5.075 80.475 5.095 ;
		LAYER M2 ;
		RECT 80.295 9.715 80.475 9.735 ;
		LAYER M3 ;
		RECT 80.295 9.715 80.475 9.735 ;
		LAYER VIA3 ;
		RECT 80.295 9.715 80.475 9.735 ;
		LAYER M1 ;
		RECT 80.295 11.350 80.475 11.745 ;
		LAYER M3 ;
		RECT 80.295 11.370 80.475 11.725 ;
		LAYER VIA3 ;
		RECT 80.295 11.370 80.475 11.725 ;
		LAYER M3 ;
		RECT 80.295 10.375 80.475 11.060 ;
		LAYER VIA3 ;
		RECT 80.295 10.375 80.475 11.060 ;
		LAYER VIA3 ;
		RECT 80.295 10.045 80.475 10.065 ;
		LAYER M3 ;
		RECT 80.295 10.045 80.475 10.065 ;
		LAYER M1 ;
		RECT 80.295 10.025 80.475 10.085 ;
		LAYER M1 ;
		RECT 80.295 12.015 80.475 12.075 ;
		LAYER M2 ;
		RECT 80.295 12.035 80.475 12.055 ;
		LAYER M3 ;
		RECT 80.295 12.035 80.475 12.055 ;
		LAYER VIA3 ;
		RECT 80.295 12.035 80.475 12.055 ;
		LAYER M2 ;
		RECT 80.295 5.075 80.475 5.095 ;
		LAYER VIA3 ;
		RECT 80.295 5.075 80.475 5.095 ;
		LAYER M1 ;
		RECT 80.295 5.385 80.475 5.445 ;
		LAYER M2 ;
		RECT 80.295 5.405 80.475 5.425 ;
		LAYER M3 ;
		RECT 80.295 5.405 80.475 5.425 ;
		LAYER VIA3 ;
		RECT 80.295 5.405 80.475 5.425 ;
		LAYER M1 ;
		RECT 80.295 6.710 80.475 7.105 ;
		LAYER M2 ;
		RECT 80.295 6.730 80.475 7.085 ;
		LAYER M3 ;
		RECT 80.295 7.725 80.475 7.745 ;
		LAYER M3 ;
		RECT 80.295 6.730 80.475 7.085 ;
		LAYER VIA3 ;
		RECT 80.295 6.730 80.475 7.085 ;
		LAYER M1 ;
		RECT 80.295 9.030 80.475 9.425 ;
		LAYER M2 ;
		RECT 80.295 9.050 80.475 9.405 ;
		LAYER M3 ;
		RECT 80.295 9.050 80.475 9.405 ;
		LAYER VIA3 ;
		RECT 80.295 9.050 80.475 9.405 ;
		LAYER M1 ;
		RECT 80.295 7.375 80.475 7.435 ;
		LAYER M3 ;
		RECT 80.295 7.395 80.475 7.415 ;
		LAYER M2 ;
		RECT 80.295 7.725 80.475 7.745 ;
		LAYER VIA3 ;
		RECT 80.295 7.725 80.475 7.745 ;
		LAYER M2 ;
		RECT 80.295 7.395 80.475 7.415 ;
		LAYER VIA3 ;
		RECT 80.295 7.395 80.475 7.415 ;
		LAYER M1 ;
		RECT 80.295 8.035 80.475 8.760 ;
		LAYER M2 ;
		RECT 80.295 8.055 80.475 8.740 ;
		LAYER M3 ;
		RECT 80.295 8.055 80.475 8.740 ;
		LAYER M1 ;
		RECT 80.295 7.705 80.475 7.765 ;
		LAYER VIA3 ;
		RECT 80.295 8.055 80.475 8.740 ;
		LAYER M2 ;
		RECT 80.295 5.735 80.475 6.420 ;
		LAYER M3 ;
		RECT 80.295 5.735 80.475 6.420 ;
		LAYER VIA3 ;
		RECT 80.295 5.735 80.475 6.420 ;
		LAYER M1 ;
		RECT 80.295 5.715 80.475 6.440 ;
		LAYER M3 ;
		RECT 80.295 14.355 80.475 14.375 ;
		LAYER M3 ;
		RECT 80.295 12.695 80.475 13.380 ;
		LAYER VIA3 ;
		RECT 80.295 12.695 80.475 13.380 ;
		LAYER VIA3 ;
		RECT 80.295 14.355 80.475 14.375 ;
		LAYER M2 ;
		RECT 80.295 14.355 80.475 14.375 ;
		LAYER M2 ;
		RECT 80.295 12.695 80.475 13.380 ;
		LAYER M3 ;
		RECT 80.295 16.010 80.475 16.365 ;
		LAYER M2 ;
		RECT 80.295 16.010 80.475 16.365 ;
		LAYER VIA3 ;
		RECT 80.295 16.010 80.475 16.365 ;
		LAYER M3 ;
		RECT 80.295 13.690 80.475 14.045 ;
		LAYER M2 ;
		RECT 80.295 13.690 80.475 14.045 ;
		LAYER VIA3 ;
		RECT 80.295 13.690 80.475 14.045 ;
		LAYER M1 ;
		RECT 80.295 13.670 80.475 14.065 ;
		LAYER M1 ;
		RECT 80.295 15.990 80.475 16.385 ;
		LAYER M1 ;
		RECT 80.295 16.655 80.475 16.715 ;
		LAYER M2 ;
		RECT 80.295 15.015 80.475 15.700 ;
		LAYER M1 ;
		RECT 80.295 14.995 80.475 15.720 ;
		LAYER M1 ;
		RECT 80.295 14.665 80.475 14.725 ;
		LAYER M2 ;
		RECT 80.295 264.875 80.475 264.895 ;
		LAYER M3 ;
		RECT 80.295 264.875 80.475 264.895 ;
		LAYER VIA3 ;
		RECT 80.295 264.875 80.475 264.895 ;
		LAYER M3 ;
		RECT 80.295 265.205 80.475 265.225 ;
		LAYER M2 ;
		RECT 80.295 221.455 80.475 222.140 ;
		LAYER M1 ;
		RECT 80.295 221.435 80.475 222.160 ;
		LAYER M3 ;
		RECT 80.295 241.675 80.475 241.695 ;
		LAYER M3 ;
		RECT 80.295 227.755 80.475 227.775 ;
		LAYER M1 ;
		RECT 80.295 227.070 80.475 227.465 ;
		LAYER M3 ;
		RECT 80.295 226.095 80.475 226.780 ;
		LAYER M3 ;
		RECT 80.295 224.770 80.475 225.125 ;
		LAYER M1 ;
		RECT 80.295 224.750 80.475 225.145 ;
		LAYER M2 ;
		RECT 80.295 223.775 80.475 224.460 ;
		LAYER M1 ;
		RECT 80.295 257.895 80.475 257.955 ;
		LAYER M2 ;
		RECT 80.295 257.915 80.475 257.935 ;
		LAYER M3 ;
		RECT 80.295 257.915 80.475 257.935 ;
		LAYER VIA3 ;
		RECT 80.295 257.915 80.475 257.935 ;
		LAYER M2 ;
		RECT 80.295 258.575 80.475 259.260 ;
		LAYER M3 ;
		RECT 80.295 260.235 80.475 260.255 ;
		LAYER VIA3 ;
		RECT 80.295 260.235 80.475 260.255 ;
		LAYER VIA3 ;
		RECT 80.295 258.575 80.475 259.260 ;
		LAYER VIA3 ;
		RECT 80.295 259.570 80.475 259.925 ;
		LAYER M2 ;
		RECT 80.295 259.570 80.475 259.925 ;
		LAYER M1 ;
		RECT 80.295 259.550 80.475 259.945 ;
		LAYER M2 ;
		RECT 80.295 260.235 80.475 260.255 ;
		LAYER M3 ;
		RECT 80.295 259.570 80.475 259.925 ;
		LAYER M1 ;
		RECT 80.295 258.225 80.475 258.285 ;
		LAYER VIA3 ;
		RECT 80.295 258.245 80.475 258.265 ;
		LAYER M2 ;
		RECT 80.295 258.245 80.475 258.265 ;
		LAYER M3 ;
		RECT 80.295 258.245 80.475 258.265 ;
		LAYER M2 ;
		RECT 80.295 260.565 80.475 260.585 ;
		LAYER M3 ;
		RECT 80.295 260.565 80.475 260.585 ;
		LAYER M1 ;
		RECT 80.295 258.555 80.475 259.280 ;
		LAYER VIA3 ;
		RECT 80.295 260.565 80.475 260.585 ;
		LAYER M2 ;
		RECT 80.295 257.250 80.475 257.605 ;
		LAYER M1 ;
		RECT 80.295 255.905 80.475 255.965 ;
		LAYER M1 ;
		RECT 80.295 254.910 80.475 255.305 ;
		LAYER M3 ;
		RECT 80.295 257.250 80.475 257.605 ;
		LAYER VIA3 ;
		RECT 80.295 257.250 80.475 257.605 ;
		LAYER VIA3 ;
		RECT 80.295 255.925 80.475 255.945 ;
		LAYER VIA3 ;
		RECT 80.295 256.255 80.475 256.940 ;
		LAYER M2 ;
		RECT 80.295 256.255 80.475 256.940 ;
		LAYER M1 ;
		RECT 80.295 256.235 80.475 256.960 ;
		LAYER M1 ;
		RECT 80.295 257.230 80.475 257.625 ;
		LAYER M3 ;
		RECT 80.295 256.255 80.475 256.940 ;
		LAYER M2 ;
		RECT 80.295 255.925 80.475 255.945 ;
		LAYER M3 ;
		RECT 80.295 255.925 80.475 255.945 ;
		LAYER M2 ;
		RECT 80.295 251.615 80.475 252.300 ;
		LAYER M2 ;
		RECT 80.295 253.605 80.475 253.625 ;
		LAYER M3 ;
		RECT 80.295 253.935 80.475 254.620 ;
		LAYER VIA3 ;
		RECT 80.295 253.935 80.475 254.620 ;
		LAYER M1 ;
		RECT 80.295 255.575 80.475 255.635 ;
		LAYER M2 ;
		RECT 80.295 254.930 80.475 255.285 ;
		LAYER M3 ;
		RECT 80.295 254.930 80.475 255.285 ;
		LAYER VIA3 ;
		RECT 80.295 254.930 80.475 255.285 ;
		LAYER M2 ;
		RECT 80.295 255.595 80.475 255.615 ;
		LAYER M3 ;
		RECT 80.295 255.595 80.475 255.615 ;
		LAYER VIA3 ;
		RECT 80.295 255.595 80.475 255.615 ;
		LAYER M3 ;
		RECT 80.295 251.615 80.475 252.300 ;
		LAYER VIA3 ;
		RECT 80.295 253.275 80.475 253.295 ;
		LAYER M3 ;
		RECT 80.295 253.605 80.475 253.625 ;
		LAYER VIA3 ;
		RECT 80.295 253.605 80.475 253.625 ;
		LAYER VIA3 ;
		RECT 80.295 252.610 80.475 252.965 ;
		LAYER VIA3 ;
		RECT 80.295 251.615 80.475 252.300 ;
		LAYER M2 ;
		RECT 80.295 253.935 80.475 254.620 ;
		LAYER M1 ;
		RECT 80.295 253.915 80.475 254.640 ;
		LAYER VIA3 ;
		RECT 80.295 265.205 80.475 265.225 ;
		LAYER M3 ;
		RECT 80.295 264.210 80.475 264.565 ;
		LAYER M2 ;
		RECT 80.295 264.210 80.475 264.565 ;
		LAYER M3 ;
		RECT 80.295 250.955 80.475 250.975 ;
		LAYER VIA3 ;
		RECT 80.295 251.285 80.475 251.305 ;
		LAYER M3 ;
		RECT 80.295 251.285 80.475 251.305 ;
		LAYER M1 ;
		RECT 80.295 251.595 80.475 252.320 ;
		LAYER VIA3 ;
		RECT 80.295 250.955 80.475 250.975 ;
		LAYER M2 ;
		RECT 80.295 261.890 80.475 262.245 ;
		LAYER VIA3 ;
		RECT 80.295 260.895 80.475 261.580 ;
		LAYER M3 ;
		RECT 80.295 261.890 80.475 262.245 ;
		LAYER VIA3 ;
		RECT 80.295 261.890 80.475 262.245 ;
		LAYER M2 ;
		RECT 80.295 262.555 80.475 262.575 ;
		LAYER M3 ;
		RECT 80.295 262.555 80.475 262.575 ;
		LAYER VIA3 ;
		RECT 80.295 262.555 80.475 262.575 ;
		LAYER VIA3 ;
		RECT 80.295 262.885 80.475 262.905 ;
		LAYER VIA3 ;
		RECT 80.295 246.645 80.475 246.665 ;
		LAYER M2 ;
		RECT 80.295 246.645 80.475 246.665 ;
		LAYER M3 ;
		RECT 80.295 246.645 80.475 246.665 ;
		LAYER VIA3 ;
		RECT 80.295 248.965 80.475 248.985 ;
		LAYER M2 ;
		RECT 80.295 249.295 80.475 249.980 ;
		LAYER M3 ;
		RECT 80.295 249.295 80.475 249.980 ;
		LAYER VIA3 ;
		RECT 80.295 249.295 80.475 249.980 ;
		LAYER M2 ;
		RECT 80.295 250.290 80.475 250.645 ;
		LAYER M3 ;
		RECT 80.295 250.290 80.475 250.645 ;
		LAYER M1 ;
		RECT 80.295 249.275 80.475 250.000 ;
		LAYER M1 ;
		RECT 80.295 247.950 80.475 248.345 ;
		LAYER VIA3 ;
		RECT 80.295 246.315 80.475 246.335 ;
		LAYER M1 ;
		RECT 80.295 250.270 80.475 250.665 ;
		LAYER VIA3 ;
		RECT 80.295 250.290 80.475 250.645 ;
		LAYER M2 ;
		RECT 80.295 246.315 80.475 246.335 ;
		LAYER M3 ;
		RECT 80.295 246.315 80.475 246.335 ;
		LAYER M1 ;
		RECT 80.295 214.475 80.475 215.200 ;
		LAYER M3 ;
		RECT 80.295 208.530 80.475 208.885 ;
		LAYER VIA3 ;
		RECT 80.295 209.525 80.475 209.545 ;
		LAYER VIA3 ;
		RECT 80.295 195.935 80.475 196.620 ;
		LAYER M3 ;
		RECT 80.295 197.925 80.475 197.945 ;
		LAYER M2 ;
		RECT 80.295 197.925 80.475 197.945 ;
		LAYER M2 ;
		RECT 80.295 195.935 80.475 196.620 ;
		LAYER M2 ;
		RECT 80.295 196.930 80.475 197.285 ;
		LAYER M1 ;
		RECT 80.295 196.910 80.475 197.305 ;
		LAYER M2 ;
		RECT 80.295 197.595 80.475 197.615 ;
		LAYER M3 ;
		RECT 80.295 197.595 80.475 197.615 ;
		LAYER VIA3 ;
		RECT 80.295 207.535 80.475 208.220 ;
		LAYER M1 ;
		RECT 80.295 207.515 80.475 208.240 ;
		LAYER VIA3 ;
		RECT 80.295 208.530 80.475 208.885 ;
		LAYER M2 ;
		RECT 80.295 208.530 80.475 208.885 ;
		LAYER M2 ;
		RECT 80.295 205.215 80.475 205.900 ;
		LAYER M3 ;
		RECT 80.295 205.215 80.475 205.900 ;
		LAYER M1 ;
		RECT 80.295 204.865 80.475 204.925 ;
		LAYER VIA3 ;
		RECT 80.295 205.215 80.475 205.900 ;
		LAYER M2 ;
		RECT 80.295 203.890 80.475 204.245 ;
		LAYER M3 ;
		RECT 80.295 203.890 80.475 204.245 ;
		LAYER VIA3 ;
		RECT 80.295 203.890 80.475 204.245 ;
		LAYER M1 ;
		RECT 80.295 203.870 80.475 204.265 ;
		LAYER M1 ;
		RECT 80.295 204.535 80.475 204.595 ;
		LAYER M2 ;
		RECT 80.295 204.555 80.475 204.575 ;
		LAYER M3 ;
		RECT 80.295 207.205 80.475 207.225 ;
		LAYER VIA3 ;
		RECT 80.295 207.205 80.475 207.225 ;
		LAYER M3 ;
		RECT 80.295 204.555 80.475 204.575 ;
		LAYER VIA3 ;
		RECT 80.295 204.555 80.475 204.575 ;
		LAYER M3 ;
		RECT 80.295 196.930 80.475 197.285 ;
		LAYER VIA3 ;
		RECT 80.295 196.930 80.475 197.285 ;
		LAYER VIA3 ;
		RECT 80.295 197.595 80.475 197.615 ;
		LAYER M1 ;
		RECT 80.295 197.575 80.475 197.635 ;
		LAYER M3 ;
		RECT 80.295 194.610 80.475 194.965 ;
		LAYER M2 ;
		RECT 80.295 194.610 80.475 194.965 ;
		LAYER M1 ;
		RECT 80.295 194.590 80.475 194.985 ;
		LAYER VIA3 ;
		RECT 80.295 193.615 80.475 194.300 ;
		LAYER M2 ;
		RECT 80.295 193.615 80.475 194.300 ;
		LAYER VIA3 ;
		RECT 80.295 193.285 80.475 193.305 ;
		LAYER VIA3 ;
		RECT 80.295 192.955 80.475 192.975 ;
		LAYER VIA3 ;
		RECT 80.295 194.610 80.475 194.965 ;
		LAYER VIA3 ;
		RECT 80.295 192.290 80.475 192.645 ;
		LAYER M1 ;
		RECT 80.295 189.950 80.475 190.345 ;
		LAYER M1 ;
		RECT 80.295 190.615 80.475 190.675 ;
		LAYER M3 ;
		RECT 80.295 191.295 80.475 191.980 ;
		LAYER M1 ;
		RECT 80.295 192.270 80.475 192.665 ;
		LAYER M2 ;
		RECT 80.295 186.325 80.475 186.345 ;
		LAYER M1 ;
		RECT 80.295 185.975 80.475 186.035 ;
		LAYER VIA3 ;
		RECT 80.295 186.655 80.475 187.340 ;
		LAYER M2 ;
		RECT 80.295 186.655 80.475 187.340 ;
		LAYER M3 ;
		RECT 80.295 186.655 80.475 187.340 ;
		LAYER VIA3 ;
		RECT 80.295 181.355 80.475 181.375 ;
		LAYER M1 ;
		RECT 80.295 181.335 80.475 181.395 ;
		LAYER VIA3 ;
		RECT 80.295 180.690 80.475 181.045 ;
		LAYER M2 ;
		RECT 80.295 179.695 80.475 180.380 ;
		LAYER VIA3 ;
		RECT 80.295 181.685 80.475 181.705 ;
		LAYER M2 ;
		RECT 80.295 181.685 80.475 181.705 ;
		LAYER M1 ;
		RECT 80.295 181.665 80.475 181.725 ;
		LAYER M2 ;
		RECT 80.295 182.015 80.475 182.700 ;
		LAYER M3 ;
		RECT 80.295 182.015 80.475 182.700 ;
		LAYER VIA3 ;
		RECT 80.295 182.015 80.475 182.700 ;
		LAYER M3 ;
		RECT 80.295 183.010 80.475 183.365 ;
		LAYER VIA3 ;
		RECT 80.295 183.010 80.475 183.365 ;
		LAYER VIA3 ;
		RECT 80.295 183.675 80.475 183.695 ;
		LAYER VIA3 ;
		RECT 80.295 184.005 80.475 184.025 ;
		LAYER M2 ;
		RECT 80.295 183.010 80.475 183.365 ;
		LAYER M2 ;
		RECT 80.295 183.675 80.475 183.695 ;
		LAYER VIA3 ;
		RECT 80.295 179.695 80.475 180.380 ;
		LAYER M3 ;
		RECT 80.295 174.740 80.475 174.760 ;
		LAYER M3 ;
		RECT 80.295 175.070 80.475 175.090 ;
		LAYER VIA3 ;
		RECT 80.295 178.700 80.475 178.725 ;
		LAYER M1 ;
		RECT 80.295 178.680 80.475 178.745 ;
		LAYER VIA3 ;
		RECT 80.295 177.710 80.475 178.390 ;
		LAYER M2 ;
		RECT 80.295 177.050 80.475 177.400 ;
		LAYER M3 ;
		RECT 80.295 181.355 80.475 181.375 ;
		LAYER M3 ;
		RECT 80.295 180.690 80.475 181.045 ;
		LAYER M2 ;
		RECT 80.295 180.690 80.475 181.045 ;
		LAYER M1 ;
		RECT 80.295 180.670 80.475 181.065 ;
		LAYER M2 ;
		RECT 80.295 181.355 80.475 181.375 ;
		LAYER M3 ;
		RECT 80.295 166.520 80.475 166.540 ;
		LAYER M3 ;
		RECT 80.295 169.160 80.475 169.810 ;
		LAYER M3 ;
		RECT 80.295 166.850 80.475 166.870 ;
		LAYER VIA3 ;
		RECT 80.295 174.080 80.475 174.100 ;
		LAYER M2 ;
		RECT 80.295 174.080 80.475 174.100 ;
		LAYER M1 ;
		RECT 80.295 172.410 80.475 173.130 ;
		LAYER M2 ;
		RECT 80.295 169.160 80.475 169.810 ;
		LAYER M3 ;
		RECT 80.295 171.440 80.475 171.460 ;
		LAYER M3 ;
		RECT 80.295 195.605 80.475 195.625 ;
		LAYER M1 ;
		RECT 80.295 195.585 80.475 195.645 ;
		LAYER VIA3 ;
		RECT 80.295 195.275 80.475 195.295 ;
		LAYER M2 ;
		RECT 80.295 195.275 80.475 195.295 ;
		LAYER VIA3 ;
		RECT 80.295 195.605 80.475 195.625 ;
		LAYER M2 ;
		RECT 80.295 195.605 80.475 195.625 ;
		LAYER M3 ;
		RECT 80.295 195.275 80.475 195.295 ;
		LAYER M1 ;
		RECT 80.295 195.255 80.475 195.315 ;
		LAYER M3 ;
		RECT 80.295 179.695 80.475 180.380 ;
		LAYER VIA3 ;
		RECT 80.295 188.315 80.475 188.335 ;
		LAYER VIA3 ;
		RECT 80.295 187.650 80.475 188.005 ;
		LAYER VIA3 ;
		RECT 80.295 184.335 80.475 185.020 ;
		LAYER M1 ;
		RECT 80.295 119.395 80.475 120.120 ;
		LAYER M2 ;
		RECT 80.295 120.410 80.475 120.765 ;
		LAYER VIA3 ;
		RECT 80.295 120.410 80.475 120.765 ;
		LAYER M3 ;
		RECT 80.295 120.410 80.475 120.765 ;
		LAYER M1 ;
		RECT 80.295 114.425 80.475 114.485 ;
		LAYER M2 ;
		RECT 80.295 116.435 80.475 116.455 ;
		LAYER VIA3 ;
		RECT 80.295 112.125 80.475 112.145 ;
		LAYER M3 ;
		RECT 80.295 112.125 80.475 112.145 ;
		LAYER M3 ;
		RECT 80.295 111.795 80.475 111.815 ;
		LAYER VIA3 ;
		RECT 80.295 113.450 80.475 113.805 ;
		LAYER M3 ;
		RECT 80.295 113.450 80.475 113.805 ;
		LAYER VIA3 ;
		RECT 80.295 112.455 80.475 113.140 ;
		LAYER M2 ;
		RECT 80.295 112.455 80.475 113.140 ;
		LAYER M3 ;
		RECT 80.295 112.455 80.475 113.140 ;
		LAYER M2 ;
		RECT 80.295 119.415 80.475 120.100 ;
		LAYER M3 ;
		RECT 80.295 119.415 80.475 120.100 ;
		LAYER M2 ;
		RECT 80.295 121.735 80.475 122.420 ;
		LAYER M3 ;
		RECT 80.295 121.735 80.475 122.420 ;
		LAYER M1 ;
		RECT 80.295 121.055 80.475 121.115 ;
		LAYER VIA3 ;
		RECT 80.295 122.730 80.475 123.085 ;
		LAYER VIA3 ;
		RECT 80.295 121.075 80.475 121.095 ;
		LAYER VIA3 ;
		RECT 80.295 121.405 80.475 121.425 ;
		LAYER M1 ;
		RECT 80.295 121.385 80.475 121.445 ;
		LAYER VIA3 ;
		RECT 80.295 77.325 80.475 77.345 ;
		LAYER M2 ;
		RECT 80.295 77.325 80.475 77.345 ;
		LAYER M1 ;
		RECT 80.295 77.305 80.475 77.365 ;
		LAYER VIA3 ;
		RECT 80.295 76.995 80.475 77.015 ;
		LAYER M3 ;
		RECT 80.295 77.325 80.475 77.345 ;
		LAYER M2 ;
		RECT 80.295 108.810 80.475 109.165 ;
		LAYER M3 ;
		RECT 80.295 108.810 80.475 109.165 ;
		LAYER M3 ;
		RECT 80.295 109.475 80.475 109.495 ;
		LAYER M3 ;
		RECT 80.295 109.805 80.475 109.825 ;
		LAYER M2 ;
		RECT 80.295 110.135 80.475 110.820 ;
		LAYER M3 ;
		RECT 80.295 110.135 80.475 110.820 ;
		LAYER M1 ;
		RECT 80.295 107.135 80.475 107.195 ;
		LAYER M3 ;
		RECT 80.295 111.130 80.475 111.485 ;
		LAYER M1 ;
		RECT 80.295 109.785 80.475 109.845 ;
		LAYER M1 ;
		RECT 80.295 126.355 80.475 127.080 ;
		LAYER VIA3 ;
		RECT 80.295 127.370 80.475 127.725 ;
		LAYER M3 ;
		RECT 80.295 128.035 80.475 128.055 ;
		LAYER M1 ;
		RECT 80.295 128.015 80.475 128.075 ;
		LAYER M2 ;
		RECT 80.295 126.375 80.475 127.060 ;
		LAYER M3 ;
		RECT 80.295 126.375 80.475 127.060 ;
		LAYER M1 ;
		RECT 80.295 128.345 80.475 128.405 ;
		LAYER VIA3 ;
		RECT 80.295 137.315 80.475 137.335 ;
		LAYER M2 ;
		RECT 80.295 137.315 80.475 137.335 ;
		LAYER M1 ;
		RECT 80.295 137.295 80.475 137.355 ;
		LAYER M3 ;
		RECT 80.295 142.265 80.475 142.945 ;
		LAYER M1 ;
		RECT 80.295 141.915 80.475 141.975 ;
		LAYER M1 ;
		RECT 80.295 139.605 80.475 139.995 ;
		LAYER M3 ;
		RECT 80.295 143.585 80.475 143.605 ;
		LAYER VIA3 ;
		RECT 80.295 143.585 80.475 143.605 ;
		LAYER M1 ;
		RECT 80.295 143.565 80.475 143.625 ;
		LAYER M1 ;
		RECT 80.295 146.130 80.475 146.190 ;
		LAYER M2 ;
		RECT 80.295 152.495 80.475 152.975 ;
		LAYER M3 ;
		RECT 80.295 152.495 80.475 152.975 ;
		LAYER VIA3 ;
		RECT 80.295 148.525 80.475 148.545 ;
		LAYER VIA3 ;
		RECT 80.295 148.150 80.475 148.215 ;
		LAYER VIA3 ;
		RECT 80.295 119.085 80.475 119.105 ;
		LAYER M2 ;
		RECT 80.295 119.085 80.475 119.105 ;
		LAYER M3 ;
		RECT 80.295 119.085 80.475 119.105 ;
		LAYER VIA3 ;
		RECT 80.295 118.755 80.475 118.775 ;
		LAYER M1 ;
		RECT 80.295 118.735 80.475 118.795 ;
		LAYER M3 ;
		RECT 80.295 118.090 80.475 118.445 ;
		LAYER VIA3 ;
		RECT 80.295 118.090 80.475 118.445 ;
		LAYER VIA3 ;
		RECT 80.295 119.415 80.475 120.100 ;
		LAYER M1 ;
		RECT 80.295 116.745 80.475 116.805 ;
		LAYER M3 ;
		RECT 80.295 116.765 80.475 116.785 ;
		LAYER M1 ;
		RECT 80.295 119.065 80.475 119.125 ;
		LAYER M2 ;
		RECT 80.295 114.445 80.475 114.465 ;
		LAYER M1 ;
		RECT 80.295 117.075 80.475 117.800 ;
		LAYER M1 ;
		RECT 80.295 116.415 80.475 116.475 ;
		LAYER VIA3 ;
		RECT 80.295 115.770 80.475 116.125 ;
		LAYER M3 ;
		RECT 80.295 114.775 80.475 115.460 ;
		LAYER VIA3 ;
		RECT 80.295 130.355 80.475 130.375 ;
		LAYER M2 ;
		RECT 80.295 130.355 80.475 130.375 ;
		LAYER M3 ;
		RECT 80.295 130.685 80.475 130.705 ;
		LAYER M1 ;
		RECT 80.295 132.985 80.475 133.045 ;
		LAYER M3 ;
		RECT 80.295 133.005 80.475 133.025 ;
		LAYER M1 ;
		RECT 80.295 134.310 80.475 134.705 ;
		LAYER M2 ;
		RECT 80.295 133.005 80.475 133.025 ;
		LAYER M3 ;
		RECT 80.295 135.325 80.475 135.345 ;
		LAYER VIA3 ;
		RECT 80.295 135.325 80.475 135.345 ;
		LAYER VIA3 ;
		RECT 80.295 129.690 80.475 130.045 ;
		LAYER M1 ;
		RECT 80.295 135.305 80.475 135.365 ;
		LAYER M1 ;
		RECT 80.295 134.975 80.475 135.035 ;
		LAYER VIA3 ;
		RECT 80.295 134.995 80.475 135.015 ;
		LAYER VIA3 ;
		RECT 80.295 137.645 80.475 137.665 ;
		LAYER VIA3 ;
		RECT 80.295 135.655 80.475 136.340 ;
		LAYER VIA3 ;
		RECT 80.295 136.650 80.475 137.005 ;
		LAYER M3 ;
		RECT 80.295 137.315 80.475 137.335 ;
		LAYER M1 ;
		RECT 80.295 133.315 80.475 134.040 ;
		LAYER M3 ;
		RECT 80.295 133.335 80.475 134.020 ;
		LAYER M2 ;
		RECT 80.295 133.335 80.475 134.020 ;
		LAYER M2 ;
		RECT 80.295 134.330 80.475 134.685 ;
		LAYER M3 ;
		RECT 80.295 134.330 80.475 134.685 ;
		LAYER VIA3 ;
		RECT 80.295 134.330 80.475 134.685 ;
		LAYER M3 ;
		RECT 80.295 125.715 80.475 125.735 ;
		LAYER M1 ;
		RECT 80.295 125.695 80.475 125.755 ;
		LAYER M3 ;
		RECT 80.295 125.050 80.475 125.405 ;
		LAYER M3 ;
		RECT 80.295 124.055 80.475 124.740 ;
		LAYER M2 ;
		RECT 80.295 125.715 80.475 125.735 ;
		LAYER M2 ;
		RECT 80.295 126.045 80.475 126.065 ;
		LAYER M3 ;
		RECT 80.295 126.045 80.475 126.065 ;
		LAYER M1 ;
		RECT 80.295 123.705 80.475 123.765 ;
		LAYER M1 ;
		RECT 80.295 126.025 80.475 126.085 ;
		LAYER M1 ;
		RECT 80.295 137.625 80.475 137.685 ;
		LAYER M1 ;
		RECT 80.295 139.275 80.475 139.335 ;
		LAYER VIA3 ;
		RECT 80.295 156.600 80.475 156.620 ;
		LAYER M3 ;
		RECT 80.295 153.975 80.475 153.995 ;
		LAYER M1 ;
		RECT 80.295 160.025 80.475 161.645 ;
		LAYER M3 ;
		RECT 80.295 162.595 80.475 162.615 ;
		LAYER VIA3 ;
		RECT 80.295 76.330 80.475 76.685 ;
		LAYER M2 ;
		RECT 80.295 76.330 80.475 76.685 ;
		LAYER M3 ;
		RECT 80.295 76.330 80.475 76.685 ;
		LAYER M3 ;
		RECT 80.295 76.995 80.475 77.015 ;
		LAYER M1 ;
		RECT 80.295 100.175 80.475 100.235 ;
		LAYER M3 ;
		RECT 80.295 99.530 80.475 99.885 ;
		LAYER VIA3 ;
		RECT 80.295 98.205 80.475 98.225 ;
		LAYER M2 ;
		RECT 80.295 98.205 80.475 98.225 ;
		LAYER M1 ;
		RECT 80.295 100.505 80.475 100.565 ;
		LAYER M2 ;
		RECT 80.295 100.525 80.475 100.545 ;
		LAYER M3 ;
		RECT 80.295 100.525 80.475 100.545 ;
		LAYER M2 ;
		RECT 80.295 100.855 80.475 101.540 ;
		LAYER M3 ;
		RECT 80.295 100.855 80.475 101.540 ;
		LAYER VIA3 ;
		RECT 80.295 77.655 80.475 78.340 ;
		LAYER M1 ;
		RECT 80.295 76.975 80.475 77.035 ;
		LAYER M2 ;
		RECT 80.295 76.995 80.475 77.015 ;
		LAYER M1 ;
		RECT 80.295 79.295 80.475 79.355 ;
		LAYER M1 ;
		RECT 80.295 79.625 80.475 79.685 ;
		LAYER M2 ;
		RECT 80.295 78.650 80.475 79.005 ;
		LAYER M3 ;
		RECT 80.295 78.650 80.475 79.005 ;
		LAYER M3 ;
		RECT 80.295 83.290 80.475 83.645 ;
		LAYER M2 ;
		RECT 80.295 100.195 80.475 100.215 ;
		LAYER VIA3 ;
		RECT 80.295 99.530 80.475 99.885 ;
		LAYER M2 ;
		RECT 80.295 99.530 80.475 99.885 ;
		LAYER M2 ;
		RECT 80.295 98.535 80.475 99.220 ;
		LAYER M3 ;
		RECT 80.295 98.535 80.475 99.220 ;
		LAYER M1 ;
		RECT 80.295 99.510 80.475 99.905 ;
		LAYER M3 ;
		RECT 80.295 100.195 80.475 100.215 ;
		LAYER M1 ;
		RECT 80.295 98.515 80.475 99.240 ;
		LAYER M3 ;
		RECT 80.295 98.205 80.475 98.225 ;
		LAYER M1 ;
		RECT 80.295 98.185 80.475 98.245 ;
		LAYER VIA3 ;
		RECT 80.295 100.195 80.475 100.215 ;
		LAYER M3 ;
		RECT 80.295 90.250 80.475 90.605 ;
		LAYER M3 ;
		RECT 80.295 89.255 80.475 89.940 ;
		LAYER VIA3 ;
		RECT 80.295 93.565 80.475 93.585 ;
		LAYER M1 ;
		RECT 80.295 93.215 80.475 93.275 ;
		LAYER M2 ;
		RECT 80.295 104.170 80.475 104.525 ;
		LAYER M2 ;
		RECT 80.295 102.515 80.475 102.535 ;
		LAYER M3 ;
		RECT 80.295 102.515 80.475 102.535 ;
		LAYER M1 ;
		RECT 80.295 102.825 80.475 102.885 ;
		LAYER M2 ;
		RECT 80.295 103.175 80.475 103.860 ;
		LAYER M1 ;
		RECT 80.295 103.155 80.475 103.880 ;
		LAYER M2 ;
		RECT 80.295 102.845 80.475 102.865 ;
		LAYER VIA3 ;
		RECT 80.295 102.845 80.475 102.865 ;
		LAYER M1 ;
		RECT 80.295 104.150 80.475 104.545 ;
		LAYER VIA3 ;
		RECT 80.295 104.170 80.475 104.525 ;
		LAYER M3 ;
		RECT 80.295 104.170 80.475 104.525 ;
		LAYER M2 ;
		RECT 80.295 101.850 80.475 102.205 ;
		LAYER M3 ;
		RECT 80.295 101.850 80.475 102.205 ;
		LAYER M1 ;
		RECT 80.295 102.495 80.475 102.555 ;
		LAYER VIA3 ;
		RECT 80.295 103.175 80.475 103.860 ;
		LAYER M3 ;
		RECT 80.295 103.175 80.475 103.860 ;
		LAYER M3 ;
		RECT 80.295 102.845 80.475 102.865 ;
		LAYER M1 ;
		RECT 80.295 105.475 80.475 106.200 ;
		LAYER M2 ;
		RECT 80.295 105.495 80.475 106.180 ;
		LAYER M3 ;
		RECT 80.295 104.835 80.475 104.855 ;
		LAYER M3 ;
		RECT 80.295 105.495 80.475 106.180 ;
		LAYER VIA3 ;
		RECT 80.295 105.495 80.475 106.180 ;
		LAYER M2 ;
		RECT 80.295 105.165 80.475 105.185 ;
		LAYER VIA3 ;
		RECT 80.295 105.165 80.475 105.185 ;
		LAYER M3 ;
		RECT 80.295 105.165 80.475 105.185 ;
		LAYER M1 ;
		RECT 80.295 105.145 80.475 105.205 ;
		LAYER M2 ;
		RECT 80.295 104.835 80.475 104.855 ;
		LAYER VIA3 ;
		RECT 80.295 104.835 80.475 104.855 ;
		LAYER M1 ;
		RECT 80.295 104.815 80.475 104.875 ;
		LAYER M1 ;
		RECT 80.295 316.555 80.475 317.690 ;
		LAYER M1 ;
		RECT 80.295 315.895 80.475 315.955 ;
		LAYER M2 ;
		RECT 80.295 315.250 80.475 315.605 ;
		LAYER M3 ;
		RECT 80.295 315.250 80.475 315.605 ;
		LAYER M3 ;
		RECT 80.295 316.575 80.475 317.690 ;
		LAYER VIA3 ;
		RECT 80.295 316.575 80.475 317.690 ;
		LAYER M3 ;
		RECT 80.295 316.245 80.475 316.265 ;
		LAYER VIA3 ;
		RECT 80.295 316.245 80.475 316.265 ;
		LAYER M1 ;
		RECT 80.295 316.225 80.475 316.285 ;
		LAYER M2 ;
		RECT 80.295 315.915 80.475 315.935 ;
		LAYER M2 ;
		RECT 80.295 316.245 80.475 316.265 ;
		LAYER M3 ;
		RECT 80.295 315.915 80.475 315.935 ;
		LAYER M1 ;
		RECT 80.295 288.055 80.475 288.115 ;
		LAYER M1 ;
		RECT 80.295 298.990 80.475 299.385 ;
		LAYER M1 ;
		RECT 80.295 271.815 80.475 271.875 ;
		LAYER M1 ;
		RECT 80.295 266.510 80.475 266.905 ;
		LAYER M1 ;
		RECT 80.295 265.515 80.475 266.240 ;
		LAYER M1 ;
		RECT 80.295 269.825 80.475 269.885 ;
		LAYER M2 ;
		RECT 80.295 271.835 80.475 271.855 ;
		LAYER M2 ;
		RECT 80.295 271.170 80.475 271.525 ;
		LAYER M1 ;
		RECT 80.295 288.385 80.475 288.445 ;
		LAYER M2 ;
		RECT 80.295 288.405 80.475 288.425 ;
		LAYER VIA3 ;
		RECT 80.295 288.735 80.475 289.420 ;
		LAYER M2 ;
		RECT 80.295 288.735 80.475 289.420 ;
		LAYER M2 ;
		RECT 80.295 290.395 80.475 290.415 ;
		LAYER M3 ;
		RECT 80.295 290.395 80.475 290.415 ;
		LAYER M2 ;
		RECT 80.295 291.055 80.475 291.740 ;
		LAYER M3 ;
		RECT 80.295 291.055 80.475 291.740 ;
		LAYER M2 ;
		RECT 80.295 290.725 80.475 290.745 ;
		LAYER M3 ;
		RECT 80.295 289.730 80.475 290.085 ;
		LAYER VIA3 ;
		RECT 80.295 289.730 80.475 290.085 ;
		LAYER M3 ;
		RECT 80.295 292.050 80.475 292.405 ;
		LAYER VIA3 ;
		RECT 80.295 292.050 80.475 292.405 ;
		LAYER M2 ;
		RECT 80.295 289.730 80.475 290.085 ;
		LAYER M2 ;
		RECT 80.295 292.050 80.475 292.405 ;
		LAYER M2 ;
		RECT 80.295 292.715 80.475 292.735 ;
		LAYER M1 ;
		RECT 80.295 297.335 80.475 297.395 ;
		LAYER M1 ;
		RECT 80.295 297.665 80.475 297.725 ;
		LAYER M2 ;
		RECT 80.295 298.015 80.475 298.700 ;
		LAYER M3 ;
		RECT 80.295 298.015 80.475 298.700 ;
		LAYER M2 ;
		RECT 80.295 272.495 80.475 273.180 ;
		LAYER M1 ;
		RECT 80.295 272.475 80.475 273.200 ;
		LAYER M2 ;
		RECT 80.295 272.165 80.475 272.185 ;
		LAYER M1 ;
		RECT 80.295 272.145 80.475 272.205 ;
		LAYER M2 ;
		RECT 80.295 274.815 80.475 275.500 ;
		LAYER M2 ;
		RECT 80.295 280.450 80.475 280.805 ;
		LAYER M3 ;
		RECT 80.295 285.755 80.475 285.775 ;
		LAYER VIA3 ;
		RECT 80.295 285.755 80.475 285.775 ;
		LAYER M2 ;
		RECT 80.295 284.095 80.475 284.780 ;
		LAYER VIA3 ;
		RECT 80.295 284.095 80.475 284.780 ;
		LAYER M3 ;
		RECT 80.295 274.815 80.475 275.500 ;
		LAYER M1 ;
		RECT 80.295 286.065 80.475 286.125 ;
		LAYER M1 ;
		RECT 80.295 285.735 80.475 285.795 ;
		LAYER M2 ;
		RECT 80.295 283.765 80.475 283.785 ;
		LAYER M3 ;
		RECT 80.295 283.765 80.475 283.785 ;
		LAYER VIA3 ;
		RECT 80.295 283.765 80.475 283.785 ;
		LAYER M1 ;
		RECT 80.295 276.785 80.475 276.845 ;
		LAYER M1 ;
		RECT 80.295 279.105 80.475 279.165 ;
		LAYER M3 ;
		RECT 80.295 279.125 80.475 279.145 ;
		LAYER M1 ;
		RECT 80.295 276.455 80.475 276.515 ;
		LAYER M2 ;
		RECT 80.295 275.810 80.475 276.165 ;
		LAYER M3 ;
		RECT 80.295 275.810 80.475 276.165 ;
		LAYER M2 ;
		RECT 80.295 276.475 80.475 276.495 ;
		LAYER M1 ;
		RECT 80.295 283.745 80.475 283.805 ;
		LAYER M2 ;
		RECT 80.295 281.115 80.475 281.135 ;
		LAYER VIA3 ;
		RECT 80.295 280.450 80.475 280.805 ;
		LAYER M3 ;
		RECT 80.295 280.450 80.475 280.805 ;
		LAYER M2 ;
		RECT 80.295 283.435 80.475 283.455 ;
		LAYER M2 ;
		RECT 80.295 281.775 80.475 282.460 ;
		LAYER M3 ;
		RECT 80.295 281.775 80.475 282.460 ;
		LAYER M2 ;
		RECT 80.295 281.445 80.475 281.465 ;
		LAYER M3 ;
		RECT 80.295 281.445 80.475 281.465 ;
		LAYER M2 ;
		RECT 80.295 278.130 80.475 278.485 ;
		LAYER M2 ;
		RECT 80.295 279.125 80.475 279.145 ;
		LAYER VIA3 ;
		RECT 80.295 279.125 80.475 279.145 ;
		LAYER VIA3 ;
		RECT 80.295 278.795 80.475 278.815 ;
		LAYER M2 ;
		RECT 80.295 279.455 80.475 280.140 ;
		LAYER M2 ;
		RECT 80.295 276.805 80.475 276.825 ;
		LAYER M3 ;
		RECT 80.295 276.805 80.475 276.825 ;
		LAYER VIA3 ;
		RECT 80.295 276.805 80.475 276.825 ;
		LAYER M1 ;
		RECT 80.295 278.110 80.475 278.505 ;
		LAYER M2 ;
		RECT 80.295 278.795 80.475 278.815 ;
		LAYER M3 ;
		RECT 80.295 278.795 80.475 278.815 ;
		LAYER M1 ;
		RECT 80.295 278.775 80.475 278.835 ;
		LAYER M1 ;
		RECT 80.295 277.115 80.475 277.840 ;
		LAYER M2 ;
		RECT 80.295 288.075 80.475 288.095 ;
		LAYER M2 ;
		RECT 80.295 287.410 80.475 287.765 ;
		LAYER M2 ;
		RECT 80.295 286.415 80.475 287.100 ;
		LAYER M3 ;
		RECT 80.295 286.415 80.475 287.100 ;
		LAYER M3 ;
		RECT 80.295 287.410 80.475 287.765 ;
		LAYER VIA3 ;
		RECT 80.295 286.415 80.475 287.100 ;
		LAYER M3 ;
		RECT 80.295 288.075 80.475 288.095 ;
		LAYER M2 ;
		RECT 80.295 286.085 80.475 286.105 ;
		LAYER M3 ;
		RECT 80.295 286.085 80.475 286.105 ;
		LAYER M2 ;
		RECT 80.295 299.010 80.475 299.365 ;
		LAYER M3 ;
		RECT 80.295 299.010 80.475 299.365 ;
		LAYER VIA3 ;
		RECT 80.295 299.010 80.475 299.365 ;
		LAYER M1 ;
		RECT 80.295 295.345 80.475 295.405 ;
		LAYER M1 ;
		RECT 80.295 295.015 80.475 295.075 ;
		LAYER M1 ;
		RECT 80.295 313.905 80.475 313.965 ;
		LAYER M3 ;
		RECT 80.295 313.925 80.475 313.945 ;
		LAYER M2 ;
		RECT 80.295 313.925 80.475 313.945 ;
		LAYER VIA3 ;
		RECT 80.295 313.925 80.475 313.945 ;
		LAYER M1 ;
		RECT 80.295 299.985 80.475 300.045 ;
		LAYER M2 ;
		RECT 80.295 300.005 80.475 300.025 ;
		LAYER VIA3 ;
		RECT 80.295 300.005 80.475 300.025 ;
		LAYER M1 ;
		RECT 80.295 299.655 80.475 299.715 ;
		LAYER M1 ;
		RECT 80.295 314.235 80.475 314.960 ;
		LAYER VIA3 ;
		RECT 80.295 314.255 80.475 314.940 ;
		LAYER M2 ;
		RECT 80.295 299.675 80.475 299.695 ;
		LAYER M3 ;
		RECT 80.295 300.005 80.475 300.025 ;
		LAYER M2 ;
		RECT 80.295 301.330 80.475 301.685 ;
		LAYER M3 ;
		RECT 80.295 301.330 80.475 301.685 ;
		LAYER M2 ;
		RECT 80.295 300.335 80.475 301.020 ;
		LAYER M3 ;
		RECT 80.295 300.335 80.475 301.020 ;
		LAYER VIA3 ;
		RECT 80.295 300.335 80.475 301.020 ;
		LAYER M1 ;
		RECT 80.295 300.315 80.475 301.040 ;
		LAYER M3 ;
		RECT 80.295 302.325 80.475 302.345 ;
		LAYER VIA3 ;
		RECT 80.295 302.325 80.475 302.345 ;
		LAYER M2 ;
		RECT 80.295 301.995 80.475 302.015 ;
		LAYER M1 ;
		RECT 80.295 301.975 80.475 302.035 ;
		LAYER M3 ;
		RECT 80.295 301.995 80.475 302.015 ;
		LAYER M2 ;
		RECT 80.295 312.930 80.475 313.285 ;
		LAYER M3 ;
		RECT 80.295 312.930 80.475 313.285 ;
		LAYER M2 ;
		RECT 80.295 311.935 80.475 312.620 ;
		LAYER M3 ;
		RECT 80.295 311.935 80.475 312.620 ;
		LAYER VIA3 ;
		RECT 80.295 312.930 80.475 313.285 ;
		LAYER M1 ;
		RECT 80.295 312.910 80.475 313.305 ;
		LAYER VIA3 ;
		RECT 80.295 311.605 80.475 311.625 ;
		LAYER M2 ;
		RECT 80.295 311.275 80.475 311.295 ;
		LAYER M3 ;
		RECT 80.295 311.275 80.475 311.295 ;
		LAYER M1 ;
		RECT 80.295 304.625 80.475 304.685 ;
		LAYER M2 ;
		RECT 80.295 303.650 80.475 304.005 ;
		LAYER M3 ;
		RECT 80.295 303.650 80.475 304.005 ;
		LAYER M1 ;
		RECT 80.295 313.575 80.475 313.635 ;
		LAYER M2 ;
		RECT 80.295 313.595 80.475 313.615 ;
		LAYER M3 ;
		RECT 80.295 313.595 80.475 313.615 ;
		LAYER VIA3 ;
		RECT 80.295 313.595 80.475 313.615 ;
		LAYER M2 ;
		RECT 80.295 314.255 80.475 314.940 ;
		LAYER M3 ;
		RECT 80.295 314.255 80.475 314.940 ;
		LAYER M1 ;
		RECT 80.295 302.305 80.475 302.365 ;
		LAYER M2 ;
		RECT 80.295 302.325 80.475 302.345 ;
		LAYER M1 ;
		RECT 80.295 302.635 80.475 303.360 ;
		LAYER M2 ;
		RECT 80.295 304.645 80.475 304.665 ;
		LAYER M2 ;
		RECT 80.295 302.655 80.475 303.340 ;
		LAYER M3 ;
		RECT 80.295 302.655 80.475 303.340 ;
		LAYER M1 ;
		RECT 80.295 303.630 80.475 304.025 ;
		LAYER M1 ;
		RECT 80.295 309.265 80.475 309.325 ;
		LAYER M2 ;
		RECT 80.295 309.615 80.475 310.300 ;
		LAYER M2 ;
		RECT 80.295 310.610 80.475 310.965 ;
		LAYER M3 ;
		RECT 80.295 310.610 80.475 310.965 ;
		LAYER M3 ;
		RECT 80.295 309.615 80.475 310.300 ;
		LAYER M1 ;
		RECT 80.295 310.590 80.475 310.985 ;
		LAYER M2 ;
		RECT 80.295 307.295 80.475 307.980 ;
		LAYER M3 ;
		RECT 80.295 307.295 80.475 307.980 ;
		LAYER M2 ;
		RECT 80.295 306.965 80.475 306.985 ;
		LAYER M1 ;
		RECT 80.295 306.945 80.475 307.005 ;
		LAYER VIA3 ;
		RECT 80.295 307.295 80.475 307.980 ;
		LAYER M1 ;
		RECT 80.295 307.275 80.475 308.000 ;
		LAYER M1 ;
		RECT 80.295 308.935 80.475 308.995 ;
		LAYER M2 ;
		RECT 80.295 308.955 80.475 308.975 ;
		LAYER M3 ;
		RECT 80.295 308.955 80.475 308.975 ;
		LAYER VIA3 ;
		RECT 80.295 308.955 80.475 308.975 ;
		LAYER VIA3 ;
		RECT 80.295 308.290 80.475 308.645 ;
		LAYER M1 ;
		RECT 80.295 304.295 80.475 304.355 ;
		LAYER M3 ;
		RECT 80.295 304.645 80.475 304.665 ;
		LAYER M3 ;
		RECT 80.295 304.975 80.475 305.660 ;
		LAYER M1 ;
		RECT 80.295 304.955 80.475 305.680 ;
		LAYER M1 ;
		RECT 80.295 306.615 80.475 306.675 ;
		LAYER VIA3 ;
		RECT 80.295 306.635 80.475 306.655 ;
		LAYER M2 ;
		RECT 80.295 306.635 80.475 306.655 ;
		LAYER M3 ;
		RECT 80.295 306.635 80.475 306.655 ;
		LAYER M2 ;
		RECT 80.295 304.315 80.475 304.335 ;
		LAYER M3 ;
		RECT 80.295 304.315 80.475 304.335 ;
		LAYER VIA3 ;
		RECT 80.295 304.315 80.475 304.335 ;
		LAYER M1 ;
		RECT 80.295 267.175 80.475 267.235 ;
		LAYER M3 ;
		RECT 80.295 246.975 80.475 247.660 ;
		LAYER M1 ;
		RECT 80.295 253.255 80.475 253.315 ;
		LAYER M1 ;
		RECT 80.295 260.545 80.475 260.605 ;
		LAYER M1 ;
		RECT 80.295 260.215 80.475 260.275 ;
		LAYER M1 ;
		RECT 80.295 262.865 80.475 262.925 ;
		LAYER M1 ;
		RECT 80.295 253.585 80.475 253.645 ;
		LAYER M2 ;
		RECT 80.295 246.975 80.475 247.660 ;
		LAYER VIA3 ;
		RECT 80.295 246.975 80.475 247.660 ;
		LAYER M1 ;
		RECT 80.295 246.625 80.475 246.685 ;
		LAYER M1 ;
		RECT 80.295 246.295 80.475 246.355 ;
		LAYER M2 ;
		RECT 80.295 243.995 80.475 244.015 ;
		LAYER M3 ;
		RECT 80.295 243.995 80.475 244.015 ;
		LAYER M1 ;
		RECT 80.295 243.975 80.475 244.035 ;
		LAYER M4 ;
		RECT 0.000 266.165 80.085 267.245 ;
		LAYER M4 ;
		RECT 0.000 268.485 80.085 269.565 ;
		LAYER M4 ;
		RECT 0.000 270.805 80.085 271.885 ;
		LAYER M4 ;
		RECT 0.000 263.845 80.085 264.925 ;
		LAYER M4 ;
		RECT 0.000 247.605 80.085 248.685 ;
		LAYER M4 ;
		RECT 0.000 252.245 80.085 253.325 ;
		LAYER M4 ;
		RECT 0.000 254.565 80.085 255.645 ;
		LAYER M4 ;
		RECT 0.000 245.285 80.085 246.365 ;
		LAYER M4 ;
		RECT 0.000 249.925 80.085 251.005 ;
		LAYER M4 ;
		RECT 0.000 256.885 80.085 257.965 ;
		LAYER M4 ;
		RECT 0.000 305.605 80.085 306.685 ;
		LAYER M4 ;
		RECT 0.000 307.925 80.085 309.005 ;
		LAYER M4 ;
		RECT 0.000 242.965 80.085 244.045 ;
		LAYER M4 ;
		RECT 0.000 240.645 80.085 241.725 ;
		LAYER M4 ;
		RECT 0.000 140.925 80.085 142.005 ;
		LAYER M1 ;
		RECT 0.000 0.000 80.295 317.690 ;
		LAYER M2 ;
		RECT 0.000 0.000 80.295 317.690 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 80.295 317.690 ;
		LAYER M4 ;
		RECT 0.000 310.245 80.085 311.325 ;
		LAYER M4 ;
		RECT 0.000 314.885 80.085 315.965 ;
		LAYER M4 ;
		RECT 0.000 1.725 80.085 2.805 ;
		LAYER M4 ;
		RECT 0.000 4.045 80.085 5.125 ;
		LAYER M4 ;
		RECT 0.000 8.685 80.085 9.765 ;
		LAYER M4 ;
		RECT 0.000 6.365 80.085 7.445 ;
		LAYER M4 ;
		RECT 0.000 312.565 80.085 313.645 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 80.475 317.690 ;
		LAYER M3 ;
		RECT 0.000 0.000 80.295 317.690 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 80.475 317.690 ;
		LAYER M4 ;
		RECT 0.000 15.645 80.085 16.725 ;
		LAYER M4 ;
		RECT 0.000 13.325 80.085 14.405 ;
		LAYER M4 ;
		RECT 0.000 11.005 80.085 12.085 ;
		LAYER M4 ;
		RECT 0.000 20.285 80.085 21.365 ;
		LAYER M4 ;
		RECT 0.000 24.925 80.085 26.005 ;
		LAYER M4 ;
		RECT 0.000 27.245 80.085 28.325 ;
		LAYER M4 ;
		RECT 0.000 29.565 80.085 30.645 ;
		LAYER M4 ;
		RECT 0.000 22.605 80.085 23.685 ;
		LAYER M4 ;
		RECT 0.000 17.965 80.085 19.045 ;
		LAYER M4 ;
		RECT 0.000 36.525 80.085 37.605 ;
		LAYER M4 ;
		RECT 0.000 38.845 80.085 39.925 ;
		LAYER M4 ;
		RECT 0.000 31.885 80.085 32.965 ;
		LAYER M4 ;
		RECT 0.000 34.205 80.085 35.285 ;
		LAYER M4 ;
		RECT 0.000 52.765 80.085 53.845 ;
		LAYER M4 ;
		RECT 0.000 57.405 80.085 58.485 ;
		LAYER M4 ;
		RECT 0.000 59.725 80.085 60.805 ;
		LAYER M4 ;
		RECT 0.000 62.045 80.085 63.125 ;
		LAYER M4 ;
		RECT 0.000 55.085 80.085 56.165 ;
		LAYER M4 ;
		RECT 0.000 45.805 80.085 46.885 ;
		LAYER M4 ;
		RECT 0.000 43.485 80.085 44.565 ;
		LAYER M4 ;
		RECT 0.000 48.125 80.085 49.205 ;
		LAYER M4 ;
		RECT 0.000 50.445 80.085 51.525 ;
		LAYER M4 ;
		RECT 0.000 41.165 80.085 42.245 ;
		LAYER M1 ;
		RECT 80.295 101.830 80.475 102.225 ;
		LAYER VIA3 ;
		RECT 80.295 79.975 80.475 80.660 ;
		LAYER VIA3 ;
		RECT 80.295 79.645 80.475 79.665 ;
		LAYER M1 ;
		RECT 80.295 80.950 80.475 81.345 ;
		LAYER M1 ;
		RECT 80.295 81.615 80.475 81.675 ;
		LAYER M1 ;
		RECT 80.295 79.955 80.475 80.680 ;
		LAYER VIA3 ;
		RECT 80.295 80.970 80.475 81.325 ;
		LAYER M2 ;
		RECT 80.295 80.970 80.475 81.325 ;
		LAYER M2 ;
		RECT 80.295 81.635 80.475 81.655 ;
		LAYER VIA3 ;
		RECT 80.295 81.635 80.475 81.655 ;
		LAYER M3 ;
		RECT 80.295 80.970 80.475 81.325 ;
		LAYER M2 ;
		RECT 80.295 94.890 80.475 95.245 ;
		LAYER M2 ;
		RECT 80.295 95.555 80.475 95.575 ;
		LAYER M3 ;
		RECT 80.295 95.555 80.475 95.575 ;
		LAYER M3 ;
		RECT 80.295 93.565 80.475 93.585 ;
		LAYER M2 ;
		RECT 80.295 82.295 80.475 82.980 ;
		LAYER M1 ;
		RECT 80.295 82.275 80.475 83.000 ;
		LAYER M1 ;
		RECT 80.295 83.935 80.475 83.995 ;
		LAYER M1 ;
		RECT 80.295 84.265 80.475 84.325 ;
		LAYER M1 ;
		RECT 80.295 100.835 80.475 101.560 ;
		LAYER M1 ;
		RECT 80.295 93.875 80.475 94.600 ;
		LAYER M2 ;
		RECT 80.295 93.895 80.475 94.580 ;
		LAYER M2 ;
		RECT 80.295 93.565 80.475 93.585 ;
		LAYER M3 ;
		RECT 80.295 93.235 80.475 93.255 ;
		LAYER M2 ;
		RECT 80.295 93.235 80.475 93.255 ;
		LAYER VIA3 ;
		RECT 80.295 90.250 80.475 90.605 ;
		LAYER M2 ;
		RECT 80.295 88.925 80.475 88.945 ;
		LAYER M1 ;
		RECT 80.295 87.910 80.475 88.305 ;
		LAYER M2 ;
		RECT 80.295 86.935 80.475 87.620 ;
		LAYER M1 ;
		RECT 80.295 86.915 80.475 87.640 ;
		LAYER VIA3 ;
		RECT 80.295 88.925 80.475 88.945 ;
		LAYER M2 ;
		RECT 80.295 96.215 80.475 96.900 ;
		LAYER M2 ;
		RECT 80.295 95.885 80.475 95.905 ;
		LAYER M3 ;
		RECT 80.295 95.885 80.475 95.905 ;
		LAYER M1 ;
		RECT 80.295 94.870 80.475 95.265 ;
		LAYER M3 ;
		RECT 80.295 94.890 80.475 95.245 ;
		LAYER M3 ;
		RECT 80.295 92.570 80.475 92.925 ;
		LAYER M3 ;
		RECT 80.295 91.575 80.475 92.260 ;
		LAYER VIA3 ;
		RECT 80.295 90.915 80.475 90.935 ;
		LAYER M2 ;
		RECT 80.295 90.250 80.475 90.605 ;
		LAYER VIA3 ;
		RECT 80.295 91.245 80.475 91.265 ;
		LAYER M2 ;
		RECT 80.295 89.255 80.475 89.940 ;
		LAYER M3 ;
		RECT 80.295 87.930 80.475 88.285 ;
		LAYER M1 ;
		RECT 80.295 88.905 80.475 88.965 ;
		LAYER VIA3 ;
		RECT 80.295 89.255 80.475 89.940 ;
		LAYER M3 ;
		RECT 80.295 88.925 80.475 88.945 ;
		LAYER M3 ;
		RECT 80.295 88.595 80.475 88.615 ;
		LAYER M2 ;
		RECT 80.295 88.595 80.475 88.615 ;
		LAYER VIA3 ;
		RECT 80.295 88.595 80.475 88.615 ;
		LAYER M1 ;
		RECT 80.295 88.575 80.475 88.635 ;
		LAYER M2 ;
		RECT 80.295 86.605 80.475 86.625 ;
		LAYER M3 ;
		RECT 80.295 86.605 80.475 86.625 ;
		LAYER M2 ;
		RECT 80.295 87.930 80.475 88.285 ;
		LAYER VIA3 ;
		RECT 80.295 86.605 80.475 86.625 ;
		LAYER VIA3 ;
		RECT 80.295 86.935 80.475 87.620 ;
		LAYER VIA3 ;
		RECT 80.295 87.930 80.475 88.285 ;
		LAYER M3 ;
		RECT 80.295 85.610 80.475 85.965 ;
		LAYER M1 ;
		RECT 80.295 84.595 80.475 85.320 ;
		LAYER VIA3 ;
		RECT 80.295 84.615 80.475 85.300 ;
		LAYER M1 ;
		RECT 80.295 85.590 80.475 85.985 ;
		LAYER M3 ;
		RECT 80.295 86.275 80.475 86.295 ;
		LAYER VIA3 ;
		RECT 80.295 86.275 80.475 86.295 ;
		LAYER M1 ;
		RECT 80.295 86.255 80.475 86.315 ;
		LAYER M2 ;
		RECT 80.295 86.275 80.475 86.295 ;
		LAYER M2 ;
		RECT 80.295 85.610 80.475 85.965 ;
		LAYER M2 ;
		RECT 80.295 81.965 80.475 81.985 ;
		LAYER VIA3 ;
		RECT 80.295 83.290 80.475 83.645 ;
		LAYER M1 ;
		RECT 80.295 83.270 80.475 83.665 ;
		LAYER M2 ;
		RECT 80.295 83.955 80.475 83.975 ;
		LAYER M2 ;
		RECT 80.295 83.290 80.475 83.645 ;
		LAYER M3 ;
		RECT 80.295 81.965 80.475 81.985 ;
		LAYER VIA3 ;
		RECT 80.295 81.965 80.475 81.985 ;
		LAYER M3 ;
		RECT 80.295 84.615 80.475 85.300 ;
		LAYER M1 ;
		RECT 80.295 120.390 80.475 120.785 ;
		LAYER M2 ;
		RECT 80.295 121.075 80.475 121.095 ;
		LAYER M1 ;
		RECT 80.295 118.070 80.475 118.465 ;
		LAYER M3 ;
		RECT 80.295 121.075 80.475 121.095 ;
		LAYER VIA3 ;
		RECT 80.295 133.005 80.475 133.025 ;
		LAYER VIA3 ;
		RECT 80.295 132.010 80.475 132.365 ;
		LAYER M1 ;
		RECT 80.295 131.990 80.475 132.385 ;
		LAYER M1 ;
		RECT 80.295 130.995 80.475 131.720 ;
		LAYER M2 ;
		RECT 80.295 132.675 80.475 132.695 ;
		LAYER M3 ;
		RECT 80.295 132.675 80.475 132.695 ;
		LAYER VIA3 ;
		RECT 80.295 132.675 80.475 132.695 ;
		LAYER M1 ;
		RECT 80.295 132.655 80.475 132.715 ;
		LAYER M1 ;
		RECT 80.295 122.710 80.475 123.105 ;
		LAYER VIA3 ;
		RECT 80.295 121.735 80.475 122.420 ;
		LAYER M1 ;
		RECT 80.295 121.715 80.475 122.440 ;
		LAYER VIA3 ;
		RECT 80.295 123.395 80.475 123.415 ;
		LAYER M3 ;
		RECT 80.295 123.395 80.475 123.415 ;
		LAYER VIA3 ;
		RECT 80.295 125.050 80.475 125.405 ;
		LAYER M2 ;
		RECT 80.295 128.695 80.475 129.380 ;
		LAYER M3 ;
		RECT 80.295 128.695 80.475 129.380 ;
		LAYER M3 ;
		RECT 80.295 127.370 80.475 127.725 ;
		LAYER VIA3 ;
		RECT 80.295 126.375 80.475 127.060 ;
		LAYER VIA3 ;
		RECT 80.295 126.045 80.475 126.065 ;
		LAYER VIA3 ;
		RECT 80.295 125.715 80.475 125.735 ;
		LAYER VIA3 ;
		RECT 80.295 130.685 80.475 130.705 ;
		LAYER M2 ;
		RECT 80.295 130.685 80.475 130.705 ;
		LAYER M3 ;
		RECT 80.295 130.355 80.475 130.375 ;
		LAYER M1 ;
		RECT 80.295 130.665 80.475 130.725 ;
		LAYER M1 ;
		RECT 80.295 130.335 80.475 130.395 ;
		LAYER M2 ;
		RECT 80.295 123.725 80.475 123.745 ;
		LAYER M3 ;
		RECT 80.295 123.725 80.475 123.745 ;
		LAYER M2 ;
		RECT 80.295 124.055 80.475 124.740 ;
		LAYER M1 ;
		RECT 80.295 124.035 80.475 124.760 ;
		LAYER M1 ;
		RECT 80.295 78.630 80.475 79.025 ;
		LAYER VIA3 ;
		RECT 80.295 78.650 80.475 79.005 ;
		LAYER VIA3 ;
		RECT 80.295 79.315 80.475 79.335 ;
		LAYER M2 ;
		RECT 80.295 79.315 80.475 79.335 ;
		LAYER M3 ;
		RECT 80.295 116.435 80.475 116.455 ;
		LAYER VIA3 ;
		RECT 80.295 116.435 80.475 116.455 ;
		LAYER M1 ;
		RECT 80.295 108.790 80.475 109.185 ;
		LAYER M1 ;
		RECT 80.295 107.795 80.475 108.520 ;
		LAYER M1 ;
		RECT 80.295 75.315 80.475 76.040 ;
		LAYER M3 ;
		RECT 80.295 75.335 80.475 76.020 ;
		LAYER M1 ;
		RECT 80.295 76.310 80.475 76.705 ;
		LAYER VIA3 ;
		RECT 80.295 116.765 80.475 116.785 ;
		LAYER VIA3 ;
		RECT 80.295 73.015 80.475 73.700 ;
		LAYER M3 ;
		RECT 80.295 68.045 80.475 68.065 ;
		LAYER M1 ;
		RECT 80.295 67.695 80.475 67.755 ;
		LAYER VIA3 ;
		RECT 80.295 67.715 80.475 67.735 ;
		LAYER M1 ;
		RECT 80.295 72.665 80.475 72.725 ;
		LAYER M1 ;
		RECT 80.295 69.350 80.475 69.745 ;
		LAYER M3 ;
		RECT 80.295 69.370 80.475 69.725 ;
		LAYER M1 ;
		RECT 80.295 72.335 80.475 72.395 ;
		LAYER M2 ;
		RECT 80.295 70.695 80.475 71.380 ;
		LAYER M3 ;
		RECT 80.295 70.695 80.475 71.380 ;
		LAYER M1 ;
		RECT 80.295 66.035 80.475 66.760 ;
		LAYER M2 ;
		RECT 80.295 65.725 80.475 65.745 ;
		LAYER M3 ;
		RECT 80.295 65.725 80.475 65.745 ;
		LAYER VIA3 ;
		RECT 80.295 65.395 80.475 65.415 ;
		LAYER M2 ;
		RECT 80.295 66.055 80.475 66.740 ;
		LAYER M3 ;
		RECT 80.295 66.055 80.475 66.740 ;
		LAYER M3 ;
		RECT 80.295 70.365 80.475 70.385 ;
		LAYER M2 ;
		RECT 80.295 70.035 80.475 70.055 ;
		LAYER M3 ;
		RECT 80.295 70.035 80.475 70.055 ;
		LAYER M2 ;
		RECT 80.295 69.370 80.475 69.725 ;
		LAYER M1 ;
		RECT 80.295 68.355 80.475 69.080 ;
		LAYER M2 ;
		RECT 80.295 68.375 80.475 69.060 ;
		LAYER M3 ;
		RECT 80.295 68.375 80.475 69.060 ;
		LAYER M2 ;
		RECT 80.295 68.045 80.475 68.065 ;
		LAYER M1 ;
		RECT 80.295 37.535 80.475 37.595 ;
		LAYER M2 ;
		RECT 80.295 42.855 80.475 43.540 ;
		LAYER M3 ;
		RECT 80.295 40.205 80.475 40.225 ;
		LAYER M3 ;
		RECT 80.295 39.875 80.475 39.895 ;
		LAYER M3 ;
		RECT 80.295 42.855 80.475 43.540 ;
		LAYER VIA3 ;
		RECT 80.295 42.855 80.475 43.540 ;
		LAYER M3 ;
		RECT 80.295 41.530 80.475 41.885 ;
		LAYER M1 ;
		RECT 80.295 42.175 80.475 42.235 ;
		LAYER M3 ;
		RECT 80.295 40.535 80.475 41.220 ;
		LAYER VIA3 ;
		RECT 80.295 40.205 80.475 40.225 ;
		LAYER VIA3 ;
		RECT 80.295 44.515 80.475 44.535 ;
		LAYER M1 ;
		RECT 80.295 44.495 80.475 44.555 ;
		LAYER M3 ;
		RECT 80.295 33.575 80.475 34.260 ;
		LAYER VIA3 ;
		RECT 80.295 35.565 80.475 35.585 ;
		LAYER VIA3 ;
		RECT 80.295 35.235 80.475 35.255 ;
		LAYER M2 ;
		RECT 80.295 44.845 80.475 44.865 ;
		LAYER M2 ;
		RECT 80.295 49.155 80.475 49.175 ;
		LAYER M1 ;
		RECT 80.295 49.135 80.475 49.195 ;
		LAYER M1 ;
		RECT 80.295 49.465 80.475 49.525 ;
		LAYER M2 ;
		RECT 80.295 48.490 80.475 48.845 ;
		LAYER M2 ;
		RECT 80.295 26.285 80.475 26.305 ;
		LAYER VIA3 ;
		RECT 80.295 56.445 80.475 56.465 ;
		LAYER M1 ;
		RECT 80.295 54.105 80.475 54.165 ;
		LAYER VIA3 ;
		RECT 80.295 51.475 80.475 51.495 ;
		LAYER VIA3 ;
		RECT 80.295 55.450 80.475 55.805 ;
		LAYER M3 ;
		RECT 80.295 55.450 80.475 55.805 ;
		LAYER M1 ;
		RECT 80.295 56.095 80.475 56.155 ;
		LAYER M3 ;
		RECT 80.295 56.445 80.475 56.465 ;
		LAYER M3 ;
		RECT 80.295 56.115 80.475 56.135 ;
		LAYER VIA3 ;
		RECT 80.295 56.115 80.475 56.135 ;
		LAYER VIA3 ;
		RECT 80.295 58.765 80.475 58.785 ;
		LAYER M1 ;
		RECT 80.295 58.415 80.475 58.475 ;
		LAYER VIA3 ;
		RECT 80.295 57.770 80.475 58.125 ;
		LAYER VIA3 ;
		RECT 80.295 63.405 80.475 63.425 ;
		LAYER M1 ;
		RECT 80.295 63.055 80.475 63.115 ;
		LAYER VIA3 ;
		RECT 80.295 61.415 80.475 62.100 ;
		LAYER M1 ;
		RECT 80.295 61.065 80.475 61.125 ;
		LAYER VIA3 ;
		RECT 80.295 63.075 80.475 63.095 ;
		LAYER M3 ;
		RECT 80.295 62.410 80.475 62.765 ;
		LAYER VIA3 ;
		RECT 80.295 185.330 80.475 185.685 ;
		LAYER VIA3 ;
		RECT 80.295 173.420 80.475 173.770 ;
		LAYER VIA3 ;
		RECT 80.295 172.430 80.475 173.110 ;
		LAYER VIA3 ;
		RECT 80.295 171.770 80.475 172.120 ;
		LAYER VIA3 ;
		RECT 80.295 75.335 80.475 76.020 ;
		LAYER M3 ;
		RECT 80.295 22.970 80.475 23.325 ;
		LAYER M3 ;
		RECT 80.295 23.635 80.475 23.655 ;
		LAYER VIA3 ;
		RECT 80.295 74.010 80.475 74.365 ;
		LAYER M3 ;
		RECT 80.295 75.005 80.475 75.025 ;
		LAYER M1 ;
		RECT 80.295 74.985 80.475 75.045 ;
		LAYER M1 ;
		RECT 80.295 70.675 80.475 71.400 ;
		LAYER M2 ;
		RECT 80.295 70.365 80.475 70.385 ;
		LAYER VIA3 ;
		RECT 80.295 70.035 80.475 70.055 ;
		LAYER VIA3 ;
		RECT 80.295 64.730 80.475 65.085 ;
		LAYER M1 ;
		RECT 80.295 71.670 80.475 72.065 ;
		LAYER M2 ;
		RECT 80.295 71.690 80.475 72.045 ;
		LAYER M3 ;
		RECT 80.295 71.690 80.475 72.045 ;
		LAYER M2 ;
		RECT 80.295 73.015 80.475 73.700 ;
		LAYER M2 ;
		RECT 80.295 23.635 80.475 23.655 ;
		LAYER M1 ;
		RECT 80.295 68.025 80.475 68.085 ;
		LAYER M2 ;
		RECT 80.295 67.715 80.475 67.735 ;
		LAYER M3 ;
		RECT 80.295 67.715 80.475 67.735 ;
		LAYER M2 ;
		RECT 80.295 63.735 80.475 64.420 ;
		LAYER M3 ;
		RECT 80.295 56.775 80.475 57.460 ;
		LAYER VIA3 ;
		RECT 80.295 56.775 80.475 57.460 ;
		LAYER M3 ;
		RECT 80.295 26.615 80.475 27.300 ;
		LAYER M1 ;
		RECT 80.295 25.270 80.475 25.665 ;
		LAYER M1 ;
		RECT 80.295 24.275 80.475 25.000 ;
		LAYER M1 ;
		RECT 80.295 23.945 80.475 24.005 ;
		LAYER M1 ;
		RECT 80.295 23.615 80.475 23.675 ;
		LAYER M3 ;
		RECT 80.295 27.610 80.475 27.965 ;
		LAYER VIA3 ;
		RECT 80.295 32.915 80.475 32.935 ;
		LAYER M2 ;
		RECT 80.295 32.915 80.475 32.935 ;
		LAYER M1 ;
		RECT 80.295 32.895 80.475 32.955 ;
		LAYER M2 ;
		RECT 80.295 50.810 80.475 51.165 ;
		LAYER M3 ;
		RECT 80.295 50.810 80.475 51.165 ;
		LAYER M1 ;
		RECT 80.295 50.790 80.475 51.185 ;
		LAYER M2 ;
		RECT 80.295 49.815 80.475 50.500 ;
		LAYER VIA3 ;
		RECT 80.295 50.810 80.475 51.165 ;
		LAYER M1 ;
		RECT 80.295 39.190 80.475 39.585 ;
		LAYER M3 ;
		RECT 80.295 39.210 80.475 39.565 ;
		LAYER M1 ;
		RECT 80.295 38.195 80.475 38.920 ;
		LAYER M1 ;
		RECT 80.295 37.865 80.475 37.925 ;
		LAYER M3 ;
		RECT 80.295 42.525 80.475 42.545 ;
		LAYER M2 ;
		RECT 80.295 49.485 80.475 49.505 ;
		LAYER M3 ;
		RECT 80.295 49.485 80.475 49.505 ;
		LAYER VIA3 ;
		RECT 80.295 49.485 80.475 49.505 ;
		LAYER M3 ;
		RECT 80.295 49.815 80.475 50.500 ;
		LAYER M1 ;
		RECT 80.295 49.795 80.475 50.520 ;
		LAYER VIA3 ;
		RECT 80.295 49.815 80.475 50.500 ;
		LAYER M1 ;
		RECT 80.295 46.815 80.475 46.875 ;
		LAYER M1 ;
		RECT 80.295 47.145 80.475 47.205 ;
		LAYER VIA3 ;
		RECT 80.295 46.170 80.475 46.525 ;
		LAYER M2 ;
		RECT 80.295 46.835 80.475 46.855 ;
		LAYER M1 ;
		RECT 80.295 267.505 80.475 267.565 ;
		LAYER M1 ;
		RECT 80.295 274.135 80.475 274.195 ;
		LAYER M1 ;
		RECT 80.295 274.465 80.475 274.525 ;
		LAYER VIA3 ;
		RECT 80.295 186.325 80.475 186.345 ;
		LAYER M1 ;
		RECT 80.295 186.305 80.475 186.365 ;
		LAYER M1 ;
		RECT 80.295 179.675 80.475 180.400 ;
		LAYER M1 ;
		RECT 80.295 174.060 80.475 174.120 ;
		LAYER M1 ;
		RECT 80.295 173.400 80.475 173.790 ;
		LAYER M2 ;
		RECT 80.295 202.895 80.475 203.580 ;
		LAYER M3 ;
		RECT 80.295 202.895 80.475 203.580 ;
		LAYER M2 ;
		RECT 80.295 216.485 80.475 216.505 ;
		LAYER VIA3 ;
		RECT 80.295 219.135 80.475 219.820 ;
		LAYER VIA3 ;
		RECT 80.295 218.805 80.475 218.825 ;
		LAYER VIA3 ;
		RECT 80.295 234.715 80.475 234.735 ;
		LAYER M2 ;
		RECT 80.295 234.715 80.475 234.735 ;
		LAYER M1 ;
		RECT 80.295 234.695 80.475 234.755 ;
		LAYER M2 ;
		RECT 80.295 234.050 80.475 234.405 ;
		LAYER M1 ;
		RECT 80.295 234.030 80.475 234.425 ;
		LAYER M1 ;
		RECT 80.295 241.655 80.475 241.715 ;
		LAYER M3 ;
		RECT 80.295 237.695 80.475 238.380 ;
		LAYER M3 ;
		RECT 80.295 237.365 80.475 237.385 ;
		LAYER M1 ;
		RECT 80.295 237.015 80.475 237.075 ;
		LAYER VIA3 ;
		RECT 80.295 231.730 80.475 232.085 ;
		LAYER M3 ;
		RECT 80.295 231.730 80.475 232.085 ;
		LAYER M1 ;
		RECT 80.295 231.710 80.475 232.105 ;
		LAYER M2 ;
		RECT 80.295 207.535 80.475 208.220 ;
		LAYER M3 ;
		RECT 80.295 207.535 80.475 208.220 ;
		LAYER M2 ;
		RECT 80.295 207.205 80.475 207.225 ;
		LAYER M2 ;
		RECT 80.295 206.875 80.475 206.895 ;
		LAYER M3 ;
		RECT 80.295 206.875 80.475 206.895 ;
		LAYER VIA3 ;
		RECT 80.295 206.875 80.475 206.895 ;
		LAYER M2 ;
		RECT 80.295 206.210 80.475 206.565 ;
		LAYER M1 ;
		RECT 80.295 208.510 80.475 208.905 ;
		LAYER M2 ;
		RECT 80.295 209.195 80.475 209.215 ;
		LAYER M3 ;
		RECT 80.295 209.195 80.475 209.215 ;
		LAYER M1 ;
		RECT 80.295 241.985 80.475 242.045 ;
		LAYER M1 ;
		RECT 80.295 242.315 80.475 243.040 ;
		LAYER M3 ;
		RECT 80.295 229.410 80.475 229.765 ;
		LAYER M3 ;
		RECT 80.295 206.210 80.475 206.565 ;
		LAYER VIA3 ;
		RECT 80.295 206.210 80.475 206.565 ;
		LAYER VIA3 ;
		RECT 80.295 209.195 80.475 209.215 ;
		LAYER M2 ;
		RECT 80.295 209.525 80.475 209.545 ;
		LAYER M1 ;
		RECT 80.295 211.495 80.475 211.555 ;
		LAYER VIA3 ;
		RECT 80.295 210.850 80.475 211.205 ;
		LAYER M1 ;
		RECT 80.295 210.830 80.475 211.225 ;
		LAYER M2 ;
		RECT 80.295 209.855 80.475 210.540 ;
		LAYER M1 ;
		RECT 80.295 209.835 80.475 210.560 ;
		LAYER M3 ;
		RECT 80.295 209.525 80.475 209.545 ;
		LAYER VIA3 ;
		RECT 80.295 211.845 80.475 211.865 ;
		LAYER M1 ;
		RECT 80.295 211.825 80.475 211.885 ;
		LAYER M1 ;
		RECT 80.295 212.155 80.475 212.880 ;
		LAYER VIA3 ;
		RECT 80.295 212.175 80.475 212.860 ;
		LAYER M2 ;
		RECT 80.295 226.095 80.475 226.780 ;
		LAYER VIA3 ;
		RECT 80.295 213.170 80.475 213.525 ;
		LAYER M1 ;
		RECT 80.295 213.150 80.475 213.545 ;
		LAYER M2 ;
		RECT 80.295 248.965 80.475 248.985 ;
		LAYER VIA3 ;
		RECT 80.295 234.050 80.475 234.405 ;
		LAYER M1 ;
		RECT 80.295 230.715 80.475 231.440 ;
		LAYER M2 ;
		RECT 80.295 193.285 80.475 193.305 ;
		LAYER M2 ;
		RECT 80.295 192.955 80.475 192.975 ;
		LAYER M2 ;
		RECT 80.295 192.290 80.475 192.645 ;
		LAYER M2 ;
		RECT 80.295 191.295 80.475 191.980 ;
		LAYER M2 ;
		RECT 80.295 190.965 80.475 190.985 ;
		LAYER M2 ;
		RECT 80.295 190.635 80.475 190.655 ;
		LAYER VIA3 ;
		RECT 80.295 190.635 80.475 190.655 ;
		LAYER M2 ;
		RECT 80.295 188.975 80.475 189.660 ;
		LAYER M2 ;
		RECT 80.295 189.970 80.475 190.325 ;
		LAYER VIA3 ;
		RECT 80.295 189.970 80.475 190.325 ;
		LAYER M1 ;
		RECT 80.295 186.635 80.475 187.360 ;
		LAYER M3 ;
		RECT 80.295 201.570 80.475 201.925 ;
		LAYER M1 ;
		RECT 80.295 201.550 80.475 201.945 ;
		LAYER M3 ;
		RECT 80.295 193.615 80.475 194.300 ;
		LAYER M1 ;
		RECT 80.295 213.815 80.475 213.875 ;
		LAYER VIA3 ;
		RECT 80.295 213.835 80.475 213.855 ;
		LAYER VIA3 ;
		RECT 80.295 214.165 80.475 214.185 ;
		LAYER M1 ;
		RECT 80.295 214.145 80.475 214.205 ;
		LAYER VIA3 ;
		RECT 80.295 216.155 80.475 216.175 ;
		LAYER M3 ;
		RECT 80.295 216.485 80.475 216.505 ;
		LAYER M3 ;
		RECT 80.295 216.815 80.475 217.500 ;
		LAYER VIA3 ;
		RECT 80.295 216.815 80.475 217.500 ;
		LAYER VIA3 ;
		RECT 80.295 216.485 80.475 216.505 ;
		LAYER M1 ;
		RECT 80.295 219.115 80.475 219.840 ;
		LAYER M2 ;
		RECT 80.295 219.135 80.475 219.820 ;
		LAYER M3 ;
		RECT 80.295 218.805 80.475 218.825 ;
		LAYER M3 ;
		RECT 80.295 218.475 80.475 218.495 ;
		LAYER VIA3 ;
		RECT 80.295 218.475 80.475 218.495 ;
		LAYER M1 ;
		RECT 80.295 226.075 80.475 226.800 ;
		LAYER M1 ;
		RECT 80.295 217.790 80.475 218.185 ;
		LAYER VIA3 ;
		RECT 80.295 217.810 80.475 218.165 ;
		LAYER VIA3 ;
		RECT 80.295 215.490 80.475 215.845 ;
		LAYER M1 ;
		RECT 80.295 216.795 80.475 217.520 ;
		LAYER M3 ;
		RECT 80.295 217.810 80.475 218.165 ;
		LAYER VIA3 ;
		RECT 80.295 224.770 80.475 225.125 ;
		LAYER M2 ;
		RECT 80.295 224.770 80.475 225.125 ;
		LAYER M2 ;
		RECT 80.295 225.765 80.475 225.785 ;
		LAYER VIA3 ;
		RECT 80.295 225.435 80.475 225.455 ;
		LAYER M2 ;
		RECT 80.295 225.435 80.475 225.455 ;
		LAYER M3 ;
		RECT 80.295 225.765 80.475 225.785 ;
		LAYER VIA3 ;
		RECT 80.295 225.765 80.475 225.785 ;
		LAYER M1 ;
		RECT 80.295 228.395 80.475 229.120 ;
		LAYER M2 ;
		RECT 80.295 228.085 80.475 228.105 ;
		LAYER M3 ;
		RECT 80.295 228.085 80.475 228.105 ;
		LAYER M1 ;
		RECT 80.295 228.065 80.475 228.125 ;
		LAYER M2 ;
		RECT 80.295 229.410 80.475 229.765 ;
		LAYER M1 ;
		RECT 80.295 227.735 80.475 227.795 ;
		LAYER M2 ;
		RECT 80.295 227.755 80.475 227.775 ;
		LAYER M2 ;
		RECT 80.295 227.090 80.475 227.445 ;
		LAYER VIA3 ;
		RECT 80.295 223.775 80.475 224.460 ;
		LAYER M3 ;
		RECT 80.295 223.115 80.475 223.135 ;
		LAYER M3 ;
		RECT 80.295 222.450 80.475 222.805 ;
		LAYER M1 ;
		RECT 80.295 223.095 80.475 223.155 ;
		LAYER VIA3 ;
		RECT 80.295 222.450 80.475 222.805 ;
		LAYER VIA3 ;
		RECT 80.295 223.115 80.475 223.135 ;
		LAYER M1 ;
		RECT 80.295 223.755 80.475 224.480 ;
		LAYER VIA3 ;
		RECT 80.295 223.445 80.475 223.465 ;
		LAYER M3 ;
		RECT 80.295 223.445 80.475 223.465 ;
		LAYER M1 ;
		RECT 80.295 223.425 80.475 223.485 ;
		LAYER M2 ;
		RECT 80.295 220.795 80.475 220.815 ;
		LAYER VIA3 ;
		RECT 80.295 220.795 80.475 220.815 ;
		LAYER M2 ;
		RECT 80.295 221.125 80.475 221.145 ;
		LAYER M3 ;
		RECT 80.295 220.795 80.475 220.815 ;
		LAYER M1 ;
		RECT 80.295 220.775 80.475 220.835 ;
		LAYER VIA3 ;
		RECT 80.295 221.125 80.475 221.145 ;
		LAYER M3 ;
		RECT 80.295 221.125 80.475 221.145 ;
		LAYER M2 ;
		RECT 80.295 248.635 80.475 248.655 ;
		LAYER M3 ;
		RECT 80.295 248.635 80.475 248.655 ;
		LAYER VIA3 ;
		RECT 80.295 248.635 80.475 248.655 ;
		LAYER M2 ;
		RECT 80.295 243.330 80.475 243.685 ;
		LAYER M2 ;
		RECT 80.295 235.045 80.475 235.065 ;
		LAYER M3 ;
		RECT 80.295 235.045 80.475 235.065 ;
		LAYER M1 ;
		RECT 80.295 235.355 80.475 236.080 ;
		LAYER M3 ;
		RECT 80.295 243.330 80.475 243.685 ;
		LAYER M1 ;
		RECT 80.295 235.025 80.475 235.085 ;
		LAYER M2 ;
		RECT 80.295 233.055 80.475 233.740 ;
		LAYER M1 ;
		RECT 80.295 233.035 80.475 233.760 ;
		LAYER VIA3 ;
		RECT 80.295 237.365 80.475 237.385 ;
		LAYER M2 ;
		RECT 80.295 236.370 80.475 236.725 ;
		LAYER M1 ;
		RECT 80.295 236.350 80.475 236.745 ;
		LAYER M2 ;
		RECT 80.295 235.375 80.475 236.060 ;
		LAYER M1 ;
		RECT 80.295 248.615 80.475 248.675 ;
		LAYER M2 ;
		RECT 80.295 247.970 80.475 248.325 ;
		LAYER M3 ;
		RECT 80.295 247.970 80.475 248.325 ;
		LAYER VIA3 ;
		RECT 80.295 247.970 80.475 248.325 ;
		LAYER M1 ;
		RECT 80.295 248.945 80.475 249.005 ;
		LAYER M3 ;
		RECT 80.295 248.965 80.475 248.985 ;
		LAYER M1 ;
		RECT 80.295 246.955 80.475 247.680 ;
		LAYER M1 ;
		RECT 80.295 245.630 80.475 246.025 ;
		LAYER M1 ;
		RECT 80.295 244.635 80.475 245.360 ;
		LAYER M1 ;
		RECT 80.295 243.310 80.475 243.705 ;
		LAYER VIA3 ;
		RECT 80.295 241.675 80.475 241.695 ;
		LAYER VIA3 ;
		RECT 80.295 241.010 80.475 241.365 ;
		LAYER VIA3 ;
		RECT 80.295 239.355 80.475 239.375 ;
		LAYER VIA3 ;
		RECT 80.295 238.690 80.475 239.045 ;
		LAYER VIA3 ;
		RECT 80.295 237.695 80.475 238.380 ;
		LAYER VIA3 ;
		RECT 80.295 240.015 80.475 240.700 ;
		LAYER M1 ;
		RECT 80.295 77.635 80.475 78.360 ;
		LAYER M2 ;
		RECT 80.295 117.095 80.475 117.780 ;
		LAYER M3 ;
		RECT 80.295 117.095 80.475 117.780 ;
		LAYER M2 ;
		RECT 80.295 118.090 80.475 118.445 ;
		LAYER M2 ;
		RECT 80.295 116.765 80.475 116.785 ;
		LAYER M2 ;
		RECT 80.295 122.730 80.475 123.085 ;
		LAYER M3 ;
		RECT 80.295 122.730 80.475 123.085 ;
		LAYER M2 ;
		RECT 80.295 123.395 80.475 123.415 ;
		LAYER M1 ;
		RECT 80.295 123.375 80.475 123.435 ;
		LAYER VIA3 ;
		RECT 80.295 124.055 80.475 124.740 ;
		LAYER VIA3 ;
		RECT 80.295 123.725 80.475 123.745 ;
		LAYER M2 ;
		RECT 80.295 125.050 80.475 125.405 ;
		LAYER M1 ;
		RECT 80.295 125.030 80.475 125.425 ;
		LAYER M2 ;
		RECT 80.295 121.405 80.475 121.425 ;
		LAYER M3 ;
		RECT 80.295 121.405 80.475 121.425 ;
		LAYER M3 ;
		RECT 80.295 131.015 80.475 131.700 ;
		LAYER M1 ;
		RECT 80.295 136.630 80.475 137.025 ;
		LAYER M2 ;
		RECT 80.295 136.650 80.475 137.005 ;
		LAYER M2 ;
		RECT 80.295 137.975 80.475 138.655 ;
		LAYER M3 ;
		RECT 80.295 137.975 80.475 138.655 ;
		LAYER M3 ;
		RECT 80.295 136.650 80.475 137.005 ;
		LAYER M2 ;
		RECT 80.295 127.370 80.475 127.725 ;
		LAYER M1 ;
		RECT 80.295 127.350 80.475 127.745 ;
		LAYER M2 ;
		RECT 80.295 128.035 80.475 128.055 ;
		LAYER VIA3 ;
		RECT 80.295 128.365 80.475 128.385 ;
		LAYER M3 ;
		RECT 80.295 128.365 80.475 128.385 ;
		LAYER VIA3 ;
		RECT 80.295 128.035 80.475 128.055 ;
		LAYER VIA3 ;
		RECT 80.295 140.285 80.475 140.965 ;
		LAYER VIA3 ;
		RECT 80.295 139.625 80.475 139.975 ;
		LAYER M2 ;
		RECT 80.295 139.625 80.475 139.975 ;
		LAYER M3 ;
		RECT 80.295 139.625 80.475 139.975 ;
		LAYER M2 ;
		RECT 80.295 118.755 80.475 118.775 ;
		LAYER M2 ;
		RECT 80.295 129.690 80.475 130.045 ;
		LAYER M2 ;
		RECT 80.295 128.365 80.475 128.385 ;
		LAYER VIA3 ;
		RECT 80.295 128.695 80.475 129.380 ;
		LAYER M2 ;
		RECT 80.295 132.010 80.475 132.365 ;
		LAYER M3 ;
		RECT 80.295 132.010 80.475 132.365 ;
		LAYER M2 ;
		RECT 80.295 131.015 80.475 131.700 ;
		LAYER VIA3 ;
		RECT 80.295 131.015 80.475 131.700 ;
		LAYER M2 ;
		RECT 80.295 135.325 80.475 135.345 ;
		LAYER M2 ;
		RECT 80.295 134.995 80.475 135.015 ;
		LAYER M3 ;
		RECT 80.295 134.995 80.475 135.015 ;
		LAYER M1 ;
		RECT 80.295 157.465 80.475 157.525 ;
		LAYER M1 ;
		RECT 80.295 149.165 80.475 151.875 ;
		LAYER M2 ;
		RECT 80.295 149.185 80.475 151.855 ;
		LAYER M3 ;
		RECT 80.295 149.185 80.475 151.855 ;
		LAYER M2 ;
		RECT 80.295 156.600 80.475 156.620 ;
		LAYER M3 ;
		RECT 80.295 156.600 80.475 156.620 ;
		LAYER M2 ;
		RECT 80.295 152.165 80.475 152.185 ;
		LAYER M1 ;
		RECT 80.295 152.145 80.475 152.205 ;
		LAYER M2 ;
		RECT 80.295 148.525 80.475 148.545 ;
		LAYER M3 ;
		RECT 80.295 148.525 80.475 148.545 ;
		LAYER M1 ;
		RECT 80.295 148.505 80.475 148.565 ;
		LAYER M2 ;
		RECT 80.295 148.855 80.475 148.875 ;
		LAYER VIA3 ;
		RECT 80.295 145.160 80.475 145.840 ;
		LAYER M2 ;
		RECT 80.295 148.150 80.475 148.215 ;
		LAYER M3 ;
		RECT 80.295 148.150 80.475 148.215 ;
		LAYER M2 ;
		RECT 80.295 145.160 80.475 145.840 ;
		LAYER M3 ;
		RECT 80.295 145.160 80.475 145.840 ;
		LAYER M1 ;
		RECT 80.295 135.635 80.475 136.360 ;
		LAYER M2 ;
		RECT 80.295 135.655 80.475 136.340 ;
		LAYER M3 ;
		RECT 80.295 135.655 80.475 136.340 ;
		LAYER M1 ;
		RECT 80.295 157.795 80.475 159.425 ;
		LAYER M2 ;
		RECT 80.295 143.915 80.475 144.850 ;
		LAYER M3 ;
		RECT 80.295 143.915 80.475 144.850 ;
		LAYER M3 ;
		RECT 80.295 118.755 80.475 118.775 ;
		LAYER M3 ;
		RECT 80.295 137.645 80.475 137.665 ;
		LAYER M3 ;
		RECT 80.295 129.690 80.475 130.045 ;
		LAYER M2 ;
		RECT 80.295 137.645 80.475 137.665 ;
		LAYER M2 ;
		RECT 80.295 143.585 80.475 143.605 ;
		LAYER VIA3 ;
		RECT 80.295 143.255 80.475 143.275 ;
		LAYER M2 ;
		RECT 80.295 139.295 80.475 139.315 ;
		LAYER VIA3 ;
		RECT 80.295 141.275 80.475 141.295 ;
		LAYER M2 ;
		RECT 80.295 143.255 80.475 143.275 ;
		LAYER M3 ;
		RECT 80.295 143.255 80.475 143.275 ;
		LAYER M4 ;
		RECT 56.840 160.850 80.085 161.230 ;
		LAYER M4 ;
		RECT 0.000 165.855 80.085 168.395 ;
		LAYER M4 ;
		RECT 0.000 173.365 80.085 174.445 ;
		LAYER M4 ;
		RECT 0.000 175.685 80.085 176.765 ;
		LAYER M4 ;
		RECT 0.000 273.125 80.085 274.205 ;
		LAYER M4 ;
		RECT 0.000 303.285 80.085 304.365 ;
		LAYER M4 ;
		RECT 0.000 261.525 80.085 262.605 ;
		LAYER M4 ;
		RECT 0.000 259.205 80.085 260.285 ;
		LAYER M4 ;
		RECT 0.000 275.445 80.085 276.525 ;
		LAYER M4 ;
		RECT 0.000 233.685 80.085 234.765 ;
		LAYER M4 ;
		RECT 0.000 231.365 80.085 232.445 ;
		LAYER M4 ;
		RECT 0.000 229.045 80.085 230.125 ;
		LAYER M4 ;
		RECT 0.000 236.005 80.085 237.085 ;
		LAYER M4 ;
		RECT 0.000 238.325 80.085 239.405 ;
		LAYER M4 ;
		RECT 0.000 277.765 80.085 278.845 ;
		LAYER M4 ;
		RECT 0.000 300.965 80.085 302.045 ;
		LAYER M4 ;
		RECT 0.000 298.645 80.085 299.725 ;
		LAYER M4 ;
		RECT 0.000 282.405 80.085 283.485 ;
		LAYER M4 ;
		RECT 0.000 280.085 80.085 281.165 ;
		LAYER M4 ;
		RECT 0.000 296.325 80.085 297.405 ;
		LAYER M4 ;
		RECT 0.000 287.045 80.085 288.125 ;
		LAYER M4 ;
		RECT 0.000 289.365 80.085 290.445 ;
		LAYER M4 ;
		RECT 0.000 284.725 80.085 285.805 ;
		LAYER M4 ;
		RECT 0.000 294.005 80.085 295.085 ;
		LAYER M4 ;
		RECT 0.000 291.685 80.085 292.765 ;
		LAYER M4 ;
		RECT 56.840 158.970 80.085 159.400 ;
		LAYER M4 ;
		RECT 0.000 182.645 80.085 183.725 ;
		LAYER M4 ;
		RECT 0.000 184.965 80.085 186.045 ;
		LAYER M4 ;
		RECT 0.000 158.970 56.840 161.230 ;
		LAYER M4 ;
		RECT 0.000 162.600 80.085 164.745 ;
		LAYER M4 ;
		RECT 0.000 178.005 80.085 179.085 ;
		LAYER M4 ;
		RECT 0.000 180.325 80.085 181.405 ;
		LAYER M4 ;
		RECT 0.000 168.725 80.085 169.805 ;
		LAYER M4 ;
		RECT 0.000 171.045 80.085 172.125 ;
		LAYER M4 ;
		RECT 54.215 153.010 80.085 153.770 ;
		LAYER M4 ;
		RECT 0.000 154.320 80.085 154.825 ;
		LAYER M4 ;
		RECT 0.000 187.285 80.085 188.365 ;
		LAYER M4 ;
		RECT 0.000 150.210 54.215 153.770 ;
		LAYER M4 ;
		RECT 0.000 203.525 80.085 204.605 ;
		LAYER M4 ;
		RECT 0.000 219.765 80.085 220.845 ;
		LAYER M4 ;
		RECT 0.000 222.085 80.085 223.165 ;
		LAYER M4 ;
		RECT 0.000 208.165 80.085 209.245 ;
		LAYER M4 ;
		RECT 0.000 205.845 80.085 206.925 ;
		LAYER M4 ;
		RECT 0.000 133.965 80.085 135.045 ;
		LAYER M4 ;
		RECT 0.000 129.325 80.085 130.405 ;
		LAYER M4 ;
		RECT 0.000 127.005 80.085 128.085 ;
		LAYER M4 ;
		RECT 0.000 124.685 80.085 125.765 ;
		LAYER M4 ;
		RECT 0.000 131.645 80.085 132.725 ;
		LAYER M4 ;
		RECT 0.000 136.285 80.085 137.365 ;
		LAYER M4 ;
		RECT 0.000 106.125 80.085 107.205 ;
		LAYER M4 ;
		RECT 0.000 103.805 80.085 104.885 ;
		LAYER M4 ;
		RECT 0.000 110.765 80.085 111.845 ;
		LAYER M4 ;
		RECT 0.000 108.445 80.085 109.525 ;
		LAYER M4 ;
		RECT 0.000 122.365 80.085 123.445 ;
		LAYER M4 ;
		RECT 0.000 73.645 80.085 74.725 ;
		LAYER M4 ;
		RECT 0.000 75.965 80.085 77.045 ;
		LAYER M4 ;
		RECT 0.000 78.285 80.085 79.365 ;
		LAYER M4 ;
		RECT 0.000 80.605 80.085 81.685 ;
		LAYER M4 ;
		RECT 0.000 66.685 80.085 67.765 ;
		LAYER M4 ;
		RECT 0.000 96.845 80.085 97.925 ;
		LAYER M4 ;
		RECT 0.000 99.165 80.085 100.245 ;
		LAYER M4 ;
		RECT 0.000 69.005 80.085 70.085 ;
		LAYER M4 ;
		RECT 0.000 71.325 80.085 72.405 ;
		LAYER M4 ;
		RECT 0.000 120.045 80.085 121.125 ;
		LAYER M4 ;
		RECT 0.000 117.725 80.085 118.805 ;
		LAYER M4 ;
		RECT 0.000 115.405 80.085 116.485 ;
		LAYER M4 ;
		RECT 0.000 113.085 80.085 114.165 ;
		LAYER M4 ;
		RECT 0.000 82.925 80.085 84.005 ;
		LAYER M4 ;
		RECT 0.000 85.245 80.085 86.325 ;
		LAYER M4 ;
		RECT 0.000 89.885 80.085 90.965 ;
		LAYER M4 ;
		RECT 0.000 92.205 80.085 93.285 ;
		LAYER M4 ;
		RECT 0.000 87.565 80.085 88.645 ;
		LAYER M3 ;
		RECT 80.295 220.130 80.475 220.485 ;
		LAYER VIA3 ;
		RECT 80.295 226.095 80.475 226.780 ;
		LAYER VIA3 ;
		RECT 80.295 221.455 80.475 222.140 ;
		LAYER M1 ;
		RECT 80.295 221.105 80.475 221.165 ;
		LAYER M3 ;
		RECT 80.295 221.455 80.475 222.140 ;
		LAYER M4 ;
		RECT 0.000 101.485 80.085 102.565 ;
		LAYER M4 ;
		RECT 0.000 143.245 80.085 144.325 ;
		LAYER M4 ;
		RECT 0.000 145.565 80.085 146.645 ;
		LAYER M4 ;
		RECT 0.000 147.885 80.085 148.965 ;
		LAYER M4 ;
		RECT 0.000 138.605 80.085 139.685 ;
		LAYER M4 ;
		RECT 0.000 94.525 80.085 95.605 ;
		LAYER M4 ;
		RECT 0.000 64.365 80.085 65.445 ;
		LAYER M4 ;
		RECT 0.000 149.345 80.085 149.905 ;
		LAYER M4 ;
		RECT 0.000 196.565 80.085 197.645 ;
		LAYER M4 ;
		RECT 0.000 194.245 80.085 195.325 ;
		LAYER M4 ;
		RECT 0.000 189.605 80.085 190.685 ;
		LAYER M4 ;
		RECT 0.000 201.205 80.085 202.285 ;
		LAYER M4 ;
		RECT 0.000 191.925 80.085 193.005 ;
		LAYER M4 ;
		RECT 0.000 198.885 80.085 199.965 ;
		LAYER M4 ;
		RECT 0.000 215.125 80.085 216.205 ;
		LAYER M4 ;
		RECT 0.000 217.445 80.085 218.525 ;
		LAYER M4 ;
		RECT 0.000 212.805 80.085 213.885 ;
		LAYER M4 ;
		RECT 0.000 210.485 80.085 211.565 ;
		LAYER M4 ;
		RECT 54.215 150.210 80.085 152.230 ;
		LAYER M4 ;
		RECT 0.000 226.725 80.085 227.805 ;
		LAYER M4 ;
		RECT 0.000 224.405 80.085 225.485 ;
	END
	# End of OBS

END TSDN28HPCPUHDB512X128M4M

END LIBRARY
